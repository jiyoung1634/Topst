PK   �z�X`)�t  M�    cirkitFile.json��_ogz���Jߙ!%�p�'{��-�ـ�$:f��E�O�|�����H���	Ĳu[�{�|qf�_����������?��O��mu���;=�����˫���i{>n�;�?.��r���������i�{�;Ο�]�ݬ����w�Ӈ�x��[����f����\.����|{��������iwx��	�����t8�<�{��&��ۯ��5ۯ�~s`�����,�j�f�5�o��>X~��W��l�f�-�c��G�o�������l��v*�d�M�_�_����ܮ����V�_�_����ܮ����֖_�_�����ޔ���������l����|ූ߭�W��l�f�-���o,���W��l�f�́uӰ�iX��+6\��s"�0��hL�V1�Ŵ��i��4�c���p�9��dv2K�rņ+6\qN�����L�j�\��W��z�a?Ӱ�)Wl�b��ĺ�i��4�i���p�9��jv5˚rņ+6\qN����M�ʦ\��W��ڦaoӰ�)Wl�b��ۡ�n�n�n���p�����f��f��\��W��\H���їҀki��4��uw3`w3`wS��pņ+�GVw7v7v7�Wl��|duw3`w3`wS��pņ+�GVw7v7v7�Wl��|duw3`w3`wS��pņ+�GVw7v7v7�Wl��|duw3`w3`wS��pņ+.�c�݌�݌�ݔ+6\�����͈�͈�M�b��8Y�݌�݌�ݔ+6\���[���P�f(p7��
����nF�nF�n���p�����f��f��\��W����nF�nF�n���p�����f��f��\��W����nF�nF�n���p�����f��f��\��W\n���������)Wl�b��#���	��	��rņ+6\q>���������)Wl�b��#���	��	��rņ+6\q>2�0�4�8�<�@�n���������)Wl�b��#���	��	��rņ+6\q>���������)Wl�b��#���	��	��rņ+6\q>���������)Wl�b���U�ݬ��YawS��pņ+�GVw7+�nV�ݔ+6\������
��v7�Wl��|duw���f��M�b��8Y�ݬ��YawS��pņ+�GG��G�H�H�I��ͪ�nV�ݬ��)Wl�b��#���v7+�n���p�����f���
��rņ+6\q>���Yaw���\��W\n�uw���f��M�b��8Y�ݬ��YcwS��pņ+�GVw7k�n��ݔ+6\�e}���������_���,J0޾����Y�?��'��8��SY��e��0y�B�S!iT:���THzPL޾��TH���<������BҨt
䩐�����<�F�� O��W��[��S!iT:��THz����<�F��L!O��o���BҨt4䩐��b�V��TH��Ӈ<��(&o%<O��Q�8��S�9a�,�
�X)O�'��;YUD��*���:�2g�:�>��1a�
}��͜Y���R#�ʹY5���73g]z'���7�ga���J�̟u靬?"�L���D+y3�֥w��x3�&}���\Z��ɢ$��tZ_���73j]z'ۓ�7�ja���J�̫u靬T"�L��AG+y3�֥w�g��Wa~-L?�Xy�
�k]z'˗�7�ka$��J�̯u�ld"�NW�u�$�]��颴>~m`~-O�Xɛ��.���Mě��0Q�c%o�׺�N:o�������_��;��D��_��>V�f~�K�d��f~-d�Xɛ��.��}Pě��0��c%o�׺�N�Do���規���_��;�5�G���<���7
1�֥w�N�x3��<}����Z��Ɏ)���Z�����7�k]z'�������}��n�tw~v����_�_3�>V�f~�K�dE�f~-��Xɛ��.���Uě��0M�c%o�׺�N�Yo�������_��;�pE��_s�>V�f~�K�d��f~-��Xɛ��.��]X�{b~-L��X�x�׺�Ndo���ت����_��;ٚE��_��>V�f~�K�d��f~-��Xɛ��.���Z��=\����:=^�=_���������0
�c%o�׺�N6qo���|�����_��;Y�E��_C�>V�f~�K�dg�f~-L��Xɛ��.��E^ě��0^�c%o�׺�N�{��ka���ʇ�2�֥w��x3�q}����Z���0���Z�����7�k]z'���7�kad��J�̯u�l#�̯�9^+y3�֥w�F�x�	�N�F܊A��>~m��Z�����7�k]z'ǈ7�ka��J�̯u�l!#�̯��`+y3�֥w���x3��}����Z��ɾ��f~-L�X9E��Z���3���Z-���7�k]z'�͈7�ka���J�̯u靬;������ywރ�����i�X^�t��SHR���g��%#�:��^��&�N�BҨt2�S!�A1	/m:�F���g�
I��Ix�@�BҨt2�S!�I1	o�TH�NF�u*$�RL�:�F���g�
I����N��Q�d�Y�B�7�Ixs@�BҨt2�S!�[�$�-�S!iT:y֩��F1	o�TH�NF�u�4'L�űc+�	�d]zg#φ�Se�\Y'Y�lY']�Ǘ5&���1����3��;y6��6�c�<V�f�K�l���f�,��Xɛ��.���gÛ)�8v�c%ofѺ��F�o&���1����K��;y6��N�c�<V�fF�K�l���fR-��Xɛy�.���gÛ��8v�c%of׺��F���*̯űc+/Ya~�K�l���f~-��Xɛ��.���g��]��銴N���k�:]��ǯ̯űc+y3�֥w6�lx3�ǎy����Z���ȳ���Z;汒7�k]zg#φ7�kq��J�̯u靍<�̯űc+y3�֥w6�lx3�ǎy����Z���ȳ���Z;汒7�k]zg#τ���Z;��F!�׺��F�o����1����_��;y6��_�c�<V�f~�K�l���v�}v��Ӎ����N�~��k#�kq��J�̯u靍<�̯űc+y3�֥w6�lx3�ǎy����Z���ȳ���Z;汒7�k]zg#φ7�kq��J�̯u靍<�̯űc+y3�֥w6�LxO̯űc+���Z���ȳ���Z;汒7�k]zg#φ7�kq��J�̯u靍<�̯űc+y3�֥w6�lx���uz�Z�ǫ��uz�Z�61�ǎy����Z���ȳ���Z;汒7�k]zg#φ7�kq��J�̯u靍<�̯űc+y3�֥w6�lx3�ǎy����Z����3�b~-��X�P\�׺��F�o����1����_��;y6��_�c�<V�f~�K�l���f~-��Xɛ��.���gÛ��8v�c%o�׺��F�o7a�iàӈ�[1�4c�ǯ��_�c�<V�f~�K�l���f~-��Xɛ��.���gÛ��8v�c%o�׺��F�o����1����_��;y&��̯űc+���_��;y6��_�c�<V�f~�K�l���f~-��Xɛ��.�����b���������x<m?-�/�?N������~��=<m����i���o����������_6�ާ�ӗ��/?>~���eW����Jok����}>�m훫\1Y�vy���u<�x��u�����2��#����W?�G(�+&��.�P��3py�b�b����ũ~�� �G(�+&k�.�P\�O=�}�G(�+&K�.�P\�O=X{�G(�+&+�.�P���zp�.�P,WL�]�x[?�`�]�X���#�<BqS?���]�X��,�<�~ o��/4�������,����Kaq�����wza�a	\n��WY�7xa�a	�n�mWY��ua�a	�n��WY��sa�a	�n�mWY�wqa�a	n���VY�7oa�a	Ln�m�VY��la�a	|n���VY��ja�a	�n�m�V� �'���@s� �>�e��[e	�Oܘ���%�>�e��[e).��W��Kx�5<�"�}�}�6,4,���-���*K�}��+4,���-�]�*K�}�+4,���-���*K�}�^+4,���-�=�*K�}�+4,���-���*K�}��*4,���-��*K�}�*4,���-���"�x���
��������k�%�>q������ٶk�%�>q�������nk���}�߿�o�wp�[������{�0а����V�,���[�0а��̶T�,���;�0а���vR�,����0а���6P�,�����0а����M�,���۞0а��̶K�,'�}�n'4�# ���vI�,�����0а���6G�,���{�0а����D�,���[�0а��̶B�,��{��{��{��{�|�������0а���6>�,�����0а����;�,���ە0а��̶9�,�����0а���v7�,�����0а���65�,W���=Ih`�n��eVY��"a�a	�n�maVY�w a�a	�n��\VY�7a�a	�n�mXVY��a�a	�n��SVY�G7�g7�7��7��7k��'�.�@�x�2ە���'n*�@�x�2ی���'�%�@�x�2ۃ���'n!�@�x�2�z,�\�wa��< ���v�,����0а���6�,�����0а������������ǧ��y{x��!ο��eq�p����Ͱ�p=�a��n��aZ���n�n����9����|ڟ/����=_�ww���'���_�����q�xx�?����~�0ݭ���f���6����a��/������r���ӧ��]z��}z�O�w��z��s��e�m^?�۫����B����w������r:>�O������p���i��fs5������Ls���fd�݌�����f����}��k7��77�qy�6���~��o�����5{�Z�`ϻ���A����x:�)��_����������+}����:������p���-ڻ�ݸ��r��OO��R����w�y7�m�k���q�a>�Űn��e����q��t�z�Z����>��}��¶�]�k����џ�|��_g_��w���B�/�����_���2����;<>��?����a�x�S���/�?8����ϻ�O��?���y����^��/
O���ߟ���?��~8�_�PK   5^�X�ZD) �, /   images/1b210ea0-4cba-494f-997a-67bd7381b5cc.png q@���PNG

   IHDR  �  
   ��.g   	pHYs  �  ��+  ��IDATx��Y�lYv��#"#�;ֽ��z"�dw�fۂ�z2 A@����2�7���O~���h�ـX$��,H���a��������7�ΰ������9��v��*�܅��q�}�^���V!��d�������>����Q��������T6?x_�_����R�V��Kyy�R�{'�k�����L�a%�.��s�B�_��W��H��Wr��Cy��ON�˅�r��ߓ��_'������̗R�{����Z�!��b#�v+�W+�t�k�x�\��+�ڵT�B|dy�X}��R,$+2=��;��w���G�ɓ'Ooct}+��J��V�?.��R���/ˇ~��k���|�\Tr���;���L�^���ޓw�粹���ǲz�J��{�����>~(��z�gr�h./��/_zt�s���=�uG~��??�X�r�V-ձ�C��r&z�'��{�s�59��ï�lq��#����\:�]'w".��Jz����ނ�����j��v)ݺ�9;}!�z&��<?{����~p"��y"��BZ�/
i�V�O_���Ǐ9oeYJ�e:������x�(��}�:��7��ן�-�l#�oWܬ/��X�[��D��A��>(>�>�r~�J6:��:9�{"�:�|���_��O�9��ח2{�D�~��'���R�W�S�>����;"�CY|U�B!�l�:�����v/�6��Ώ�|���^�Zx�z�~�����}?�-��?��TU%y��~������o�������v-X��C����3�yt_l6<d>��ڎ�>��NV:w��5�����=��V
���[ouݗ���-��e�{m#A?ۻ�\63���̗oIY�x�A�=�#�g���8ރ�6?����ڲ}������ʂ��Ϲ�����U�=;�Ϲ�p|f}y!���4Mõy||�y����0��o���܎O5n���h���?�:��ʃ;�2S ݜ}(�j-��3y�$t�� `��Gw�J��y:ݔy)Ǉ��� Tt3�f���!�*��	l4|D��`�"V
��ذ��]hhp���s�9���x ���-s��*P ��Eč�o8?�/	���}��CX�xN����H�2W���~��ù���"�"Վ����'��o{���������F�����5F!��C��ۀ��^� }��p%���Q��U��q�\�g��r�0x�ñ�ǝ������A&�g|#�3�{q�2��k��sN���Rx���c(8;���K��> ���(�x�[�s�ysQ1�x��^2�����Bns�����7��S�ec:g�ޛ 5/S�y�@�ӥ��lͧ��=��JM��w�?�����:��?��e���3$̦kٽ��#��S:O����L�����s8=����'r;>��޿�qy���W���=~|(��������{.^-�Eu(-�F��V��^�0��T!��s%��B�%4hz�ZFj�@�ݨ���f�%##�͚��ͥ�O �jн
���sjv������ZO iW[*l�A ��e�R���37XY�h0�{i�'k#m�\Xn	�񝖚�����P��b���w{�� 	��P�v�mUY�AB �}/�;iڍ�
��n%G}�7��h���$���ތ0 �]3,�v�J��gv��_�nV|?�-�
ez�f��R����iL��k����
�ڵ�pv��Z��M�,W��"ǿ{����ϖpL�ͩ��Ϫ��I熥����٩��tWz�-��w�ST��[����=y�����H���?<�t�O0~�3*Qi�<�W|��.ikY|�b�B�h��T>��|ʍ��������Ǥ�j�zg|�)]�Y�Q��ܿ�7�E��;Sz�͡O�h��M��l\�!�àH�fΦ����������x�
������?��_�7Y������T:�tW�^��s� 3�4.U��K7���[�"pU^fR�����n"�f� ��W`\oL*�t�����n������3Y��fk]
M!��e!����X���M���m�(p�V�-��X.� i.Cb,����`�%P�{�6��\��=8�[Uxx��J\�L:����h�{XQ�Zi�`��\��+��@��:k۵�m-��J��R����J ,g�Q5��<����p?����K�.U�9�ȅ�^�B�7��yf6?�%,|1�c6���6oi�l��X�x�_S�D��]�^WJZ��j�z<��>�֫�c� �̯@�չ��<-V��n^+�+o��q�d{]��Z���:�H)�8W2��-���a�t��J� �wH���:��ν����1 ��o&
�3e�̓#�+z�
-]ߺ�U����}�����(�3�@L�^{o�s�ֆ�s>����I�;Ql�����M�MR؆W\c�=t��x��4[��k�W�"�܎O=n���`���O���}��R���+i���Rv�r�`&�6D[�wT�������B6>�E} ����A���V��-A�Q��i:�GP ��*`�¬3�6_��������V��J��
�w�n���R��{)�*\�t�[;G^u
��M�6>,^�?#w ���c��:��<#���[��,
4�,7��C���# CI�ĥśsn�=���|X�y֪�\Jޮd���f܌�Ly��E.I`��#��~..��9_���KY�_H]�%�8���g�\r-�ş��E��U�b�	xoR\nz�����X81�efJ ��9��\�|:��<*v��ߩ¢+�n� L����^�ܦQ��t�w��p��r͌�#�-S��G�QM��d�����}o:�V����y��`"�!�A1`�f�OTvt����ĵ���G��uo�$0��{�_�����$��%DOKTp�I&#@�c���MZsܗ1���tQ!IJ�����J�����<����-�~����?��y����ɱ�n�֪
�#pjm��9]�V"��ey����%��-k	x)�����K�@:nX~@��8�� |+�nUt��P9�,�H���7H�k�*���%[`���'n�`1�m4h�d���bUi�'�MsUVkV�_���Jc/��fR�jC�+/��!x�{ \��S��\�TQ����C�U)���ʖB�7 �m�V����<x��S0hl�6Y镛�W�z���
��l.�y��]D�N���$���Bu"��q���7�/_�`2;&	%���|{(y>��7����P�=�kz,��B��u���_����8�K�7��|Uq�sؘe���F��^�d;-H�]�F�2L�����@+>M��b���|������2rCX�e�v��gVP�ɣ�ʵIP� ���"s�>=�x9����2Dn��T7?���8��x=��z��;Ƃe F��~�s��t;ּ�␾G�Y����\&�ZR�����������x?��G�����fu�['�A�5���]^����\7��z��/$S�Y̜�N����]̥�*9z�m��H1W�Wz�(�Ȃ��V���T,,}E��7�"�j��3�H	U��i�1�����HڏMb$�1�� ,0$�*�:�X'ܘ���C�S8t���j�0���Z'��E���r�<���,̃�C'�y��.ޠ@�:��mĲ��u�e��h}�h������,���/��n٢4V.��$��� c��s�4b�s������fN��b!HZY��c����R�0�k�Z]f�_�t{���9U�2�7��� <��/�lp���$4��H��5<7<%b�s�'�M�j��D��u�&��[#�A��iz�	��D?�<��N�a#�� �b�y�/z_�yBLˆp ��c�u�P|4�+����y�|�DP X]&{��kŋ�׸�1�:h0�o����I���roƥEt$Kf>=�����Y�I����U�;��^��r;���x?�q�������Z���s	땬��%��R��x� � P�*7�88�l����S�7ɋ�wrW.�/�Wj	�����B3݅��3�w�UfD��48��"�;1g�;q�p���(�I���8�4�I�
{\��� Z�!�s�k( ����gnssW{�,ܥbn|e�v�%׹+��Zt1
��r����)���,^lbHL�%��"۱�p�� � ��lq?����W>�w]vtW���kVΞ��?\Di�'{��9���WAQ�DA��P�\�ђW%��������ʘ�EQ9z=�lMw5��T�H}�5���?��fׯu�R�� ��~����g5�/�/�a�\:xY�����@x�q���z�������#/ �D� ��u=َ�[9IN�j5a����ɄY|ߏ3�uj�����'���U���T�a�v_��g�x v��fJ�������9h������~��{G��k6�jpm$4�Z$NfK9<<��公t�Vj���'�ߝ�"�y:��;^ʬ�����g��L(��_��\�wT��$?��i&ܠ[�5��.��9����rrS���})'''�!�S�C^���/G�Cc�Fw3����1��� ���g�Ϛ,���@��Zj��B�l#��HU�\�x�w��J#Je��\�G�r��0������ܨ��-�?��:���h'��ݞ��)��T �˄�1�!�R'n`(3��D��y����<LY"0G�E!օ�d��	�_��0w�8o��BK�G�2�f�rs��b���uk�s38�R�P�e��B���Gg	�:�`-�rS��G!�U����'Z�x���^�=lާ�ӂ�^Kon�)�&�����ߘ+��cϪ�<�\� ���N��ES`ٷ��:�2�'�p���wpnd������Kم��Z��ߊJH"QaE�G�k�~,@��<����|aJ��O퉀ۇh�N%�.H�k[���f��<R��m�􇘒�� M|��֫=�i�(}'��4O�}OU,�O������9���}m�����\W��"i�ѥV�
� L!� )6
�ܗ��wa�u�$��-6�
J�g;��h5@V���\�b.5	29ٮ.�8��ЇхeZ�~�Qd���ؒ��b�>�[R�Uj����l&xFݕ �N���}_h�;�gq�dy{1+V&-�HD٢H�5 �g�E�:<��L�LM�����"ݵ�|��R�md�[��,	,��6Ę��]w %����a�4z� �9�ͬ^2s�(�h�g�>2ݳJ?S���B9�g�����"����Do
 Ĭ(��C�yȂL��ٰƦ�̜	�� ��(�p1$��r�c1�&)�Ļ��-����������Z��h��x-�Z�X/~�Z��k�����W� �{�8/���#H|�Q$��%�p6<�t-��K�`��g������R��17�;0e�O�������-~|�q;q��x�죿S�ݪ�-�z<GΧ
�y9#����Th\��r��"e��S��~�*\,�Л��Í���-�]��&���s����=�!���q.���r�v��IN	�<\Z���a�n6�5�=Gf����(���!���k`�t��6jE���A�G	V�GM8=�Z1|C@����DW�4����
�hy&�H�rcd	dm^��f���s��k�rTf�Xi��%[�h�n�����R�ma�G� t̎D1]G�r����MB�8ޤ^#�:g�W�S���4��p�+����x���s"�
.غ�Wo�`����;�P�?ߴS:xޥ�E+8�;��cD`��m�Q��C̅���<"VE�ւ�[�!��S�AQj,���\Vt��u�l�L�x_~ �1�d�u��Uܫ���V��t�����ݰn��2"�k?���KIڷ�/=n��s�����?������=Y��۲�J�!���M:�-e~x,n����JZ�/�o�ݡ�i�;�~���kd�!���}�G�N�蒬�\D�X}"L�(�������t�����TU�\�P����&榍�3�"$�/��-���8i���"�
sk��٬��{D)IT�
H��%��U'.
�N��"`�2ˢ���b��`��D&\ʴ/�$����ps�����=�)�W�OcR~�D��R���	*w-���s6=�k�3��)!��I��y9P(1L0�BL�2���y���B1 �EУ�W�7%Ez����U%	q^�TIq���]���a�Qa�R]�F��j^�/yt�:?�x�4v����"�a�����ЍM�CDR��V��ᘞ�|�Ve���9�Tp�c�@dЧ��zq��&A�.1�(q �>�����M�ȝ*������T!N�;e�O~wY������9��?��o]]]|��iͥ��Z6WW$o,e����"�R���K1_�:��ڈ,zT�xuK�k��7��{�6���i\��S7�1�s�֍U��&A��5�@{���l��쳣�j�0����q�r��t��ե���[Z�ƺ�r�f1��c=�n� ��a~,e�'��,�q��+B�Ә�`�F�,M.Xn�&UK���L%���q�dd$�h��2�Xe�̘l��*��>
��-x���& I��[PB��b��8�>Vc��E�[���B�n!]�<CbJG����Ұ:@7�+}�Uj=G+��eZ틇�6y�֚��X�
i(������*/��1�=�[�ʒ�aN�4�����t�n�M�<�}�,�t'���E����q��qp���+]+��՛���+i�FK����`F�s���lO���F}!nP�$�TPA·���p�� ��,��6�g�|�7x���4�~��t\��@tj������Rfa!�����C�
�
p;cm��6)j�2�K��h�
�h~ W� |CFk��-G���!X;F��Ga~?ʑ,mh۬y=��1�$b婮�M�c����}�9��e�c���E�s�Z_2Eh��ڣ2Va��Ab�	�O��ݨ�RA�!.	#H,�������ͩ.� R���Ǻ՘K��]+�-�0VVb�I�����rbǸ���0��2Wݴ�"]�Vd��L	]��<�N���t���'`=��IGf�>����`�ǒ��ü����Q�C�*y�����
Lpo���k��#*}�r�k^����d�^�7��DW�44q�~R��V;[�)���Vu��7�c�s�]�J��4#=����2�ޯTѸ��ޘ/J�]b���۵B���4�_�z���&���]��1\��O�ۿϝ�W7 �b���O9n��s�����?����gGR*����G�5�.�Y>�yv rt$��T��n���9��܇*�rnd�.�	L�v`M�fqX����$8��*����9�GY�l�25A3�U|I,�+�@��OE3�֝U��w�V!�ɲK%��N��X�z#m���X�#Ty򋽑���fC��r����c.h�ՋlHV���y���M�yC�	�;�[
{g��u�=b`}YL�B�ET7
�$��^��N�MނQ������F7�]�g����D�>1��9s*$�`� �,^#_Ų\��EnR�2Z/���5��ݐ:��c���F�^&�"�����ąlkh��L�"=�O:nrO�]&�H!��vc��w= �K�{���1��}��~(��U,�m�2U	;i�,�E��3������ي�H�Js�]�')XC��-��y�im�)m����<�*ݩ�<��nǧ���9��_�tݷ�ɼʥ��|O�~[˝�5Ax�칥ͨ�TW�+P`e�C<-X�7J����2��XJU�Y�*��rs3��裻ld؎�zV2]��ݻ�[�?	ƴ�`F �Z	S��w5�[H�Y����+2Z��$��6^�1�յ@�Q�F4���6d���Uf��huV�>�p^�y�g�H=Z3;���\�.��p��n#֘[�3u	���f�Dj�Z��o���y{�؉�퀳g��=�ȼ��yk)&S���K���4�����d������PlqK4��kT�ye1�mI�����DK|���k�*/%� �h1hA󽹹٥����<0"��mI��ԝ�:kw�X�wA�O��s�A(,p5o��;�X�C$*AF�L�!p����s��[��o�NS]�Kٻ~Rxi�k��Ʊ_�]���;>���a��'?��:o�/Pf����|.�Z���(E�_I�j��y��90����_X��4 :�l�fL�#�@`�N�e�rΎyHet#S�*`!���OpI�C.)��5~����������
p}״	ˢ�����>�3�R��Vlr}�]lNZ��F���Z���r��ݷ���)�\
����B����P��*���\����&Vk��y��*�ql䆆)#HYY[��܊[@�o��D�f�Xo=+����L�<H��1�<����Moi1�Z��������88r!k�cn�j!�"�ϥ�f�Y�.����2m��a�sjM[��J�5�*�;�bVb��O�`���y�\��~�䑀����y�]E�� xt��e����n#(M�z�\L2Ů���&����Vx+qjgk����|(݈
\�����eb���G��"�W��OA?Y�3*^]���G�潈�����ݳs�,�/�٤#�~�*�]�,�us��?eN�1_8VKc��R̚�;z�B�ۜ����s�`x�b�]g���G~Z�"�L�h���5��l��<X{߅��Tɟ�%��&�[o�_v���0�_<��G(���.�RC�[䟗Ym)8�b�-�tS44��2�c����r%�\b�j7��J�b?��B�[�ԛ�QŘ�D��S�P&�ߥ��Κ'@a��gΆ�5k1'�)�o����ߍq�������?�� �2���[���p5W�ׄ(P�`f�MU� "��V�f�'�ܬ@&HQ�0����\�����{}���5��:V|Y��sJ�ق�t�t�5�c߼��nA�x�j�G��Ůi0f���M���.q �
,0���Y�c���Bj�%F���_0�%ճv�r�%��&�&��T����4��{JjJĭa���*b7��p�7xƿ������T |�|�N�,�D�I� #����݀���϶6��X2�xuт����1!�O�F\������M]����}��4B����U���ǧ����}�{������o|���x�f���M @��5t�!������QX�h7Iհ�t�1tS)GhĽ�BBx���YGل�S�p�iԘ�1ʯ`,���bC�)�b���מ9�԰c���:n_��D���07*�IzC*̞�����
h ��5��S��i2�����M&yMQ(������cz�>E{=z�_;�\4��~(ݗ�S�E-ʱ(�56���'������b���)+nQ��㓳���V�Yk����-��q�
������b���ɤB�/��x�k>��Hl���^�~��޼|�s^S��M��v�J�&�##{S��'����`t��ld�?��x�t����0��S�w���m��)����+텽XpE��?*{z�u}k�~�q����\\|���;�|v��H@As�y%�nL�zk�V�n�b�r��3+����ʭ�?���^�E�� �U�VsxWe���l�p�c��|t��՝ط9.��������1�v�Ɵ2�{�>��ػ6D��\C���P^3R6
���Q����_6�Q`��IG%��:
E���<�齄(�ܞp�cm�)9�������U��L O��t;�'K��
M	��*bp�pS\=�%�k#�=�B��>����4?%�g��#�cO�n��c�i�v�1�H"��Y��dO�����c9B��%��\����U����L����M����χ�7���O*��1�a�yZ�D_c��s�s�����t�^�CcV��9�P�Ɗa�z����'AN�붮��	����T�,�v|�q����n�����|@(]>��6
��a&m����F��s�.�Y�����\"V��@�w�Oy��Z��/�blae�c�T`$��Ʌ̈\�l5y�|s��!�j�|Okfbd�T�
��,�wр ��ɪ�nc����jbA�|L���3�{:t�qc�I��>ѱ���a�n5� ���Er��X�/���@�:�Hz7Y���4G9��`ꂟ  a��ޜޏ.�!�]��u2��KPvAdd��c�X؃���^�d]؝`�b<(�[�ɔ�˜o�� ��H��#*0��G��G�r���d��tPdT8XeIv�,2�m}��>�~�q���^���?��'��6�Z��\�nC�7������;��e��[�{�3z:��H������f��>Ĭ'�2�{S♂n���Pnǧ�����������?�ÿ}rt �
�YU�f}�#!p�{	�ޑ>su%��~[i�6,�F��`��Q�)S���B��U�B7!��T�����pE Ixi:�%�6�7�"�.�BB����v~�qͭ�Y H�æ�˛��t��
8�6vv,��k�^���t\�G��*P"��|enyƅ57�V���s���ߧ�\,@��=�����=�2XnM0̽k��Y���.y*�m=�3��5�3^w�$ w-���]�v�~�c�g/�.���������l"tnǋbϒwY�ce3;WR ���ڊ ���-�C�3�9�z�q�L�g�X�I���3v.�s�}�ݏS�d�?�ܙ�>���q�R����9�j���Λ����׷�ܹ>�sfi�V%���U]�)��������!��+�Uzߏ�v|�q���X����~���b^JUf2�+9�ZQ ����l)��6HZ�$l�v#�R摹(B�uN3����k����~Ip�C��7�Ջ�	�۩�٪���R�(}Ԡ�]+�bM��;���כ��% IqY�1�Y�nI�4,��DkS�X���,a���,(����S*z�@���]]��67�5	A{dLg���z*��{
$.r��/6s�'@�,���Ra¬(�z��b��@A��z�.1����\�!��Y�1E)�o��~L׍�O ��@�*�5ZPk8r�&�R���e5��|��v�,ΰLߘzn�O�͏D�Aaz�;v',�1�`G����{��\����A���ց�|Y�t��5�@��{�ȥ:㙑���t����H'�-�����k��}b����3^o7rp`l����-�v|�q���h��� �v^�B��Q��jzYΎX��`VK�Z���iZ+c,��:�=ja�z��*2MC^�ېVlKЅ�:1�1��1�XL.�]H�|U{�#K%����By�I�ٮ[*սM�&xj�L9b� WZ���K�hue�o�5n�5����[�\X�LyaI͖��|7/���]̄�K� �(Xu/�Af���<\L��=����T@a(̊�%�2L	Vx�$�E�2�a�%n����ט����������x�	�X���5F���Ec����N���=>���V�X�It�F0�fY�] H�1����u㓂hz֟��6}N����Rgs�	 �eV!-��p���k��]w���i|썜1-.�����@���%�1-�q㥻�����(�^^^��|���ޗ���-�~������&,������<��}Z�}�,�E��~�f?R
9��Pa����@-�b���ཚ�b��� �c�`�*�|EY�G����\�5� vG�x.�I��E,`���%�a��c<L`�Tl��x��SOީ�v�הץ�߮7����I�G�ޢ�klz+$K���Uk�T�"|[X��e����e���\бS����Z}z��]��}�����_�7l#����w��s���td1m������z~ϟ�X����%��q�<Z󇇇rzz�s����čl������/ǚ��e��q6��j}�a�M@ͼ��- ~���W]ȶ�V;�I��C�x�Y�N\�=ױw�x�np��5���T39}v_!<�si�� }o����L��C-h�A����f�wK0�0n����<��: !�v���s��G��+��bf���i6\��a}sC$a"u��.Ow1!��GO�����[�f�"l�֏\H�2[����`�'/���u�z�����S�}���p>��/��������*�혎[�������4�lkj����w@�'6��lby?����&���µ�R�k�5i��/�sf�Yޣ�F�uhśz����l�A ��d �4��"��b���֫�s�J)�]r��Ҋ0n�����9��.cU-]WPf�87�����G�f�?�.g^/�S{?�I�JW��Fw*���|Nu���o��|��7Z����Tz ���\��b -�S���9�7��[b�������غ���C@�Z"�؍�Umf�,w `�\㻬�7>�4�a���-��a��fݝww�}_�����@�us<e,"�C*��� �R�b$�ųX���\Ê]�[��7�=�T�#^B0F���P���/��9=s�'��݉'�u�]���\���� ȍ����@�:�O8X��ط���w�}���������ޒ�,��4����Re����<5�QnLG�pQ�lH�<�p�Z(a����P#�"+Y��q��>zs ��*X�ʹ�rBA�*A`��A)���U\,"`�R�2$�)ob5'c�y3��0���\V�LfX�
WT�_�Z��i��JN"���HC���a��'�*ݼ.k���&�:��7�s;F�.>���5�@%���&�L��#N�ݔͽ?�'K�����M�ki*����V�ʢ�.�s���,c�8of ��O�y� ��3�ԯ,9 ӹ�O�{��������z���z���ߦ�M�d�V��len�x��xby��PQ�?�:�Є#����	a�Mo���kt�ο�=c�!�?�`��X���.�U�K�l|���2��"�C���@����0��x��1׺��V�n&����?���O_�]��W��]�,����������xsuU���Oʫ��Le������}��_�_���_�{����Y��y����ί�}G7�Z..V�P��S��z)��R,4����j�Ϋ����c+	�����A lM��>E�
HI�)�����1'6u�E�Z0� ��{ ?��T�纋xje�.��7�|ɲm��[�슔ǎ+V�����9���iU�akno��������#��,	���c�㵍`����Y��Q��1���|Qs���5%���X۴n�5������� ���X�{�-m�4��}(��[Rb�Ìe��$��J�+���u�����1�z��~��2B���z� @)N|���m7����~�u�=�"���X��G���D�PaMפ��Ř�\m7��C��}��}��"�ey��C[No
�_/��o��㞺ؓ+/0���O;(�v0���_?^���|��>��o�����˳Ws�A�Bŀ��{ǇGrp|,GG��\����ӟ���_��W��|��-�~F������ݬ]k�BsĠk�Z�bq"\ƨ6�ca���e� ��j�V3���JZ xt3��5�QEP�d�m����y#&1^'2�{g��3�����ݬZV��˙^��<븺����V�~�����{&�v�%L@}Լi�;"��J � ���5�1�l$�Y	N+ZO��X���I(�>qg"�I����`�e�Ś/�������s�/X�up���`9�Q��r�o��n�n;�5<GoW���ļ�,(L$�`�+��c�3���=������v�YhX�,*_.�ڊ�$e��P�blt���=�����{�
~���5�����YO���b�QS,YJt�s<�&z��w��1�}�A�s�Y�>l��j1����]�Pכ���,h�YpL�{���IU���X�`�u �e�܃��Rِ�Ҏ^���q��j7������o��w���/..~����߶}���V�Fl{y������\�<y"��淢gñ���_����s��s���7s��g0�����ڦnļԅ��%�%T���=q��Z�Ř%�G��F�ٜ*� S�utp,a�$��v]n ��t��(,}���U��u�W�p)='���jZ� ��7���d*�޲=b��q�\�n���՜�e���7�Fk �0��p�2`m,a���ͦX% �7"ON�z���N��b�;�&��B���ҽH�!� 6_ ��:$���K�Cb�_�Nu��®!)5�$,�X�$tiR�*�Z���F!ZȆF�c���6z6z�Iaֽ�\�����=�9Fr������	�
b���B��6O�+ιKka���Hm,�����Ua��r`]���{�����ޛ�O�En,��,����ڒ���x��z;k|߫"���r����K����e]˽���q��{�~�^����Y���ف�O�{�kʊ��/�����|�s�.��i��0��]�O?���z�Y�w~�w�׾�<��j��Lb�3��*���+U�U!��ϟ}����������[������ɏ���S�QZ�d�.�i���]�MQZ��ꃁKZ�M�Y]��w���o)�b��n�}͘\��+�BI��rf�fY4� M�\�T���w��
hL~ڨI�X'�!�����+�ǝ���h	�x�"a��X/�=�B�3�f,��+�
C�9���rM�}��d�(�c	�7�,�&F*��y6�B0�g�88�j�[�V~3Υ��+SKdwN���Hk)g�#��a�kXD0�b�3Q�T9c���sL�B��,6����J�[��3������)cyd��Ks�g/��lt�d�&V3��
������`�U�&w�x�$�˓��|���u��t�;Z�E�f#��ZvkU^;rl�d�K��5�\���|��c�=���(���� �3������>%D���5�����LHs���p%�Wۿ���L�z�H�z򘹾���ʡ����^���s����v�B�N�Q�Լ��|x||�e�����g\��������2�.��V�a���b��낋�9�h.�
"��ق,h,\��%���n�j�Z�!V��
�3i�Z�ٚ��u����Lx���[A	�\]�ѧƍ�z��I��.9�j�BnR�x�`ta���w4�<��3�c���lm���;+~����J�ˢ�4�.�߬�tc����q����ΑZ#hq'-7>�!�OW�b����0������Va��<:��;G2/f��E]��%�����X� �	ҽ︺o�#7VѺ	���8kt"$(@�g����M^<W�s���i��(�lTAlt}p��*���Έ�S�uF��:��]@̞��X���g������D:�f3z<��
��}O�cl;)�����J�B(e6���We֯��h����A͇�Ƙ>�s�!	�I�����z&9M�T����X:g����A*� z:jc吘��@�쩄8�Ӎב���&??*=V��H��z���!�]�9�K /-]���G/ �V_/_������3y�w��q�CpU�2F|lWct��*�2�8�z��m�G����2n��������e���n�E��u^}��_?w����Y�����i~xPK���<9���_]JUߓ@�� ��
� �f��Y�ҝ��Z@��h�<XXE�0D���9PaU�wd%K}o�r���/#/�Ś����^��܏����e��B�I��R5�颷�Y���m���
�FϿޮ�������L-�/^���٩�U�Fd���U�ȣ���bG��;+�A0��7D����%�����D�@,���L�p���lVHK����J�����r���n�J7.^�C.G�w�nk���0*�Ԧ� �-��Pe6H;�)n	�-�f�y-w�:f���
�9-�����N�j1K�VbQ!���d�%�0�"V.���>ݶ�3 ^UZ1{a��{(+�S|�tz�HdFB3K�	߷��F��νZh,�󗣒��3��K���l����S-$BU�y�3X���5�eO����zlAq`����m�mQY( �k�{�H�'K�;\��i��+$zߔ:6��-5�H���3y*'��#��V�?X�bs�9V0D��E�d�8<O9V�
���ͽ��[�SP���,#,��b˚7P t�*ۂ�E�>���NO'0�ّ,�we�Ұ��.�R�<�����l�uʬ�dP����x�g\<���0e�k$�>��3�B1!����>븆*������F� '@ؿ��ҏ�@l׺W��}�r���\��A���۬;]��\��QV������?�X�u]�Q�c��������;Ϟ={���g����������O~z�4M�w���xy��?�������?�颞��ѝ�?9::z����/E~�h����T@���������<y|��՚c�e8%�nf4��t�e �����fU�ڥ{����w��RnT αq���>�X����B!��TAILxy���E��27u���5��$6׎1I�GQ��C�l���ۇ�Xg[�ut�Yk�n�|����v��	l>S�TT�g.�5\�pX�p���l6+���*��`�ѩ��s2�]l kW�Ҩp@7�P]��?��%}�V\�Q���a�,j��x����ev��T`�h�"x���Xu�X����h0_���V�r�r!6O.�T�/����w�&/(�'�77k� ����Z<�y�1]��,����X��U���ױ
X#��3ٮ�lW�Q&CJ�S�Rk���YUW��8γ��V��ޗ!���i�k��rx|�y��J�չ<X2�1�]�	~?��&E��rK��h��<a��"ѽ�����zR�ӻ�|d�%�'��o
�*�WD"���@�}2��}=�����T�f�չR�9�����sN��]��.|T�C���f�,��*B�b�ԥY��}�^�~�3�_�׼^���"8i�<�0ײo��(��4�gs�3��7�r�`�w���0���NNN�(����|
�^�q�[ȁ{U���.Pw&���W�4n�7���{����_����Y�����|�׿�����p�����]^\|.G,������Ç�o?yr��/}������o����v��o7탾i�%�fdk���c���m�T���٪�Pm/ߨ&�fx��Oi*�2Z�&��
5�2�UH�Y��C]�(0�#���[P��6m�T��)
A.���{q?�JTQ3}���r4�K�	;��li#D��s��qF#�X�)����Ft��*�=ko^�&��D�u_�g�3���e��3����N�J�YXx�j���lQD7}Nwn�Vҭ^ɺY��qA�u�Z�:0^ς���b\�LƘ,�`.g J �ؤ���t���1�B�.��]'��9DE����!6Eǋs�EJh�c�h��%��0@��e}lZ�r�do;Z�����`6� Y	VNf�c�3�d�b�A�U�ox�K��Z�=-dc��wsq����Ρ�-+�J��ɍ�:���W�)g?� �D�2N���z�5Z�%yE]o5*��6_8������X���deJU������ѵ �*x��D� ٷ�pqΦ�������.˭��=�;v^*�P�A,�˲�:�P�g�R�2�
U�@fbl\���W��4��0q����j�:�
dm)/_^J{�y��~yx,�y�����\�o��LZ^}nզ���x�1d� S!�HWp}�0�I�cw4���ŅZ�+���k
jlT�\����z������</�[��y�˓C��<���>�R/7�Q�P�P��>?}yO�k�Ea6�oW��������oȗ����w����?�3y��9�B��T9_,����{�'�`A~gu�fIB�Dl6k��TS�.`q:�l�>,��B�n�z��l���f3�a%E66h�7z՜䂂2g�H��
�Rf�%]�I��i�XP�3d�BXw�b��/a���.�,7��g+����&0�=},o�c���?�P�9���	C\���tT�������c|�����e���*2!�+�R�.��-]���
�j�����gR�� ��""��M�Bߋ�.��% �h-���-p�,����,��FP},Dw�3y�Ɔ�|�Yڸ�V�g*]8�w�e�Rk{u �����bn��Q[~.�����B8FV�3V��t.rX>�h�g)�`�D�Z@�
��
h}uT �{)W[U��L� 
7�TA'�-�C�����r鐶ӛ���Y�Txuo��:��A+\����Jf��,����Z�.Z�zd����2�u��jt�Q���K�w�7N?�x����`��a�b��T�n����<��2�
 B)�`��D��F��f���3(-�*P>��n�#��j�ry��y�f'��i��*�..������\"�G\E�S�����KNHa��`���2�>b
P g�4�Лp��TUk�����g�չܮ:�ەʱ?�����?��Ϟ���\��?x�}IZ�K�]`�#E
mG�xa]O�3=a(�S����Ν;�ч����
֙|�-�
A�����?����<<>�61A�:����_�u�ַ�Z�Z�-�Ie����֭|�W�N��F7D���r��='�'$@VY�F�>�d���J7��k��+�V5�M0�a2��ݮh� +�Y�U ��Y4��`��7���Ӎ�|9�cO]��z۬I:��&���\�U�k|�x�grx�d���ѡ<|x_�˥ԋ"��X�QJ�����n7p����h��9��Ď�a�C[F�ټ�YAk����F���T�.�3k��z��Vn���K�R�V�3�Xb2Dpѹ��*P�M^I�h��#�/��Cn�|�Ѩu�La���u�r�A%��-���ղ �ި.Wİ؆ ���xYo��O7<�՘��p�5��:0�9��1s�=�P�ݞ.P70�	� W�zɈM���p��݃�},�阳]&2 ��0���pU�p�<�t�{��c/Ȋ�y���&����>ӗ�͟����PG�;\���K�A٫О-I�c�HUR�j^�~��تeu��XP��=X�.�z^,j�ݑ{�Q�K��i������::l宜(�TT��������(�_P���g�k���K�WTb���z�#��:#ށ�公T!���&�p��\��L��ٕZ���:��i���
f^�*)]WKS���݈��e��9^�3���<���p=�������9���z����t���..X�UNE|���n�՝�V5�E0D�5�����LI���Ȱ��^���ַ8�/_���?���]��y٪ppx �AU+d�5�b�+�9��_φ���Go�7���B�p��U���Қ.��e��G?���o=|�6�|�"�����V�ri�^�
s�0�Bְ��z�D�o?6_�E�ۉ0�1ݮ[I{y)Ŧg�e�lD-�E�p�����L�P�� �k��(/"�Q�S��(Z�W�Õ��6kY�=��顥뷶4���fYoT�����Nŧn�\7�9��R�M2�-��kU���C�P��ѿ�i-�� Xo�C�0�V-M��l����Q�dw:\�}���v�W w�*l������97pj�9M|��G{�̫ ?�ׅ��g�/ղ�U���c�sF��:9�x�\����G
���[�ִPKw�X��W��T�����:��g^�xF�������x�>���c�`y](0,�zQ3���%~�k�R-���\+0��~V��R
2<��,�Q�"\��y0F,�1���WϞK��e�j��0.n�3���ϥu[��;��ܟ��Y�i�O�|���%�A,�H�m˸�wֱ����\��
`S�L�&㔬>c��������*2ꭂ�%���lG�oF��lq@��u��+���OP����U��3*/kX���N�?�����D!mo6��3�����"���%�O>ӥ>7 /b�t�K hᳫ��{��������V�ST)��:�-d�u�dW$�!ݍ�8��q�'�QWT��t�Ō��V����~Sn����\1��<��!z���6zƜkO�w	�`D|`�l�-$l͐�H��3�Db.�5��w�$��k�����CC 1Z�����G1�ö�$�.zi�G5\����~G�ݿK߶��ޕ/��^��z�+q��{��jytB�ݬg
��Z�.Xdh��\u�.��j�`�>{���.6�Z=z�d!���4��GE�~� ���Pa_���`�`S�$$�g*`50'B��f� %��&�#֌�*�l��j	�`i�dիM�˙j��EM�cI�@����K�k��2ּm�!o�Z������i�������7��9�
h��O������&E2܍ ��x�8t0!�Y�$|���_�o�*�Ҭ�n��ѳ�����\d��
3�9N?~!A����W$W��WR��Z���ՙ���]�Bt����X�0h�t�JN�η�Rm�輫����V����g���<�8�M��^��ϗ$����9?�P`\�.?:��8;Y��\�����%�y��nu��@��]�u����{�� �x����3�P`���v||O�yM�K╂��Wr���jsE�~���g	�[�0�Y�V�^1b�-\,m< �V�No�?\J?�g������x�Uӊ�FfwU��Wz���\���u�:��U���H�Q]a���~%S�d9�
�7�΂Q\��F+<�y�p�@aA!�d�a���|����F��^/,<�/�\�P$�
�{�ui�c�eq���1.��0�xqb�����Ŀ���K�֦����ʱ"�B���ʭ[齫�K`�0F��U�Uk�82GV1��|�m?�7���c
��sQ���Tx3��eH$p�3,,׽��uJ9��I�U��^\��!���V�!���÷�׾��rtrl���8W���@)�z>ȎTU�x =d�Jgx2�܎����������[��>3Chpp%S�)Ђ$Qͬ��ܕ�i �,�v�Y���{���p�`�ߑt�
��[2=4>��
��
1��@��I�j� 5�)7H��U�&T�X)K�O��� d�Z@
f�n���䳒q�m�+�6�P�h�c*k��/.����@�;�"�qkvO����GjM���5곗�r�X�B-���=��j��1:W$AA��s���r�V`V+�J7�Ďޚ4* �������g��?�Sn4� 1�stL���1��)HܻwG��,X�R��|([�^_�P>�4����]��/.i�a|�`Z�z^�S��*;��
��E�x��C}>����E�Lq>W�U�z�Q�~��=�� ��ř��s*Q��5S���K�)�
����JM�z����@�c�YG<OT�B�p�5=[��
��B���>�vh@��^��{r�U�4�1�B5��sY�ta��-��)*8_��e��`n(�>���?s�_5+�P��zSk
�8���(����k{���ȮP����b�P���Fe8�@�Q�
u���:�&��t0����B"���@���.XkE$���Դ\�zk����`���n.�v1S�X��|�k%/DL�³�,�j��"��
L-,P�R�����TC�������k�ΰ?;~�,b�1q�=��4ʂ�V9�&�B�]-#Y�(ˡ(�X��
�Ы�R�k�X�'c��Y�Ӵ�,fbd���" ��D������C�����P(���mUY���M�.��F�M�j{�O승]G�5�d����,����=W��f+��T(�,G��(��GG����"aI���Z(����a:@��ɭ:P1?����Q����],Ok5��q���q��ၬ+
��*=�l������Z���e�t����x֍��j�:��])�]����F�v-sy������B��G
|,%��r��߹j��~��rt�D�A�;���Fz��5�)�Uy�ّU�0��� 	d�����ogО-�7#���;_Q �R�`^�`.�Q�|�7$ �/aي�zI�bA��y�p�����ѫ�]x&� Ή�6�_z��?=Ν�``*x�����V7��I	dY��q3+���t���b�)����T��CxQ ��s?�)L�D.6@��g��>����������xK��rx�mk~�Rcu��V-�v��uf�tF��4n�TƖs �需��y�s�{�b�����r� �YS�?T�bqv�YD�)I�G�M�g��VcS1RZ���+�M����r�9��4�$�$*�n������To?����'�ئ����t%h��Ŕg�{J�2,d6�ք��-�]���b�Og9��7�#��X�wk�;k�i5�q,4I���ʲ!�,s�Td�)�
2X�R��������ٯT��N����(֬%��qM�-�Flp��Kz�����||��Liĺ�Po��u)�}��է&�kPl�8<�3]�d�����CX1��ˡE�V5�#�`6��-7�d�6��U��[��t��_����K�=:Q�R�3���Ժ��t���s��+���cY�w�(�yg0����8�6��7�=���Ͷ+��L|��_��1�{���>��Z�Y( �'��ά0b�jA>z�15WT((| ��L��ͽc9T�ɓGL%b~l-�h���,��RD8c��*�S�ϯܙ��@xp|"3U"hyVH�4�8��:�8+4Y�L,?؛����<Ƒ�b�4$�����2D{>���4X���B	 �Y�-��`�����t���2��*_�� ���B- �X�8Re��b0��	�T��H,�`��`�+�I�1�8 ��*<��v~��Z٤l'-C-ӗ�k�fݱ68Sk
G ���|A���d#���9<N6(0����M��x��	��,N�Z`�Vj,�#6�K1�gt6����RaJ�7�`�a��s�O��{�#�P�	V�i�����Y,�b�w�����c����#U{@���j�����9�l(�[�+�P�-����|����l�\�1m�U�����i7��~F���8��>3~'e%L�;�&K#ȱWv�IV��'��uB�k�'e4���������|A�-������γ�/dvth�1�RA�B�Z�R�d���a!j��j	\��d��/�>�_|�\^�z!��o�U[RS��㇏��[O���̲7n�2��-�+ٰzY��s�}$��tM�,\�[��6�!��V�9�l5{��:�呂|�Y� ���(L�@�`C2�_�����o(�7�ۛ���E*�3K�בR\��!��`��F�)%�L�88�W.d���FnbyC2,��b���8�~�(A��Ҏ��U�Xd@l�"��c��R;�zK�#�0Άkh(׭"�s�B	IY�̾A��0�uˣ��b����&��E�4�h=E7'b�I��w4g͇�c�P���[�2�Pyb ��͆EGR���9+\�[wx��1ň���b�
�UY��N�bg%��c�`Ƃ�9�vl����!]c�|�r���Z�G�jrg���&����tf���E�@a5��\�����3�w
t���+�d�0*u�#0����c��%9'��Y��:]T���!]�=_.K=��z�c���kZ�:^߀���c���o��`����e8��}*=?���l}Ht]g{U:�����9����zS�S^�$N�œ����\��g$���s*M�k�P� ��}�у�����|���-w�')��]Z(m÷�Ea\�/�+�W��G_�����'��r��£�O���{����R,e���w�{|pG��<��kղ��FM<U7�X���������X�fA�1�Lq���ji��e��Y�����EWg����rg��� ��v�D]G����ZSBj�g)/)?����+P��*30�n�h�ٞ�I`)N�;O��ʳJ\�I� ���"�,����X�Y�V����5�}�����0ܗ��ɀ�n��Bv@��ǜU�9�Hھ��b��@�� �=S)tp�Ȕ��' ���N,�AX�<���0�����KE�w-6+#ʪ�$2y��᥀ MSFK����c,q��"��ެB���hi��Y���)�|*K<�2��/��X'��䱿�wC.hzM�����Y�c�����1VkeGk<~��yJTvĔ�8aT�XC+,�1_o�A��m�u�_h%U�ۿ��j|�{8��ܛ�W�d�b�~ҩ{S�1ݲ0σr���s�w[^�4�rc�3M�����/<�^n6����������#�]nZ8p1�߃�]U=I(���j��ta~�����z�W���[�<^ʼ��V����&�Dr��	z $t�n*����ds�;D+)��C���?0>!�f�c�tc��)$� �Hވ��#�NMۺ�xg�/c���FI,.�+����iS��Il	 ʦ���0Ū3���w�Բ!�F���&��3�yq��F��Z(�L�{K�]��X#~,Q����m������@K��ZI]�t����V�D��su�~��K�.ZF�5�'��x/�Q�ܲo��ľ�1�^��w6�����]a7���t��,��g��2�ǷL�1�΍�K��,]j`���!�\���M��k�E�=#=��q�`�������"?*Cq	�e*��;�_N��}P�w{�`!�{�H��Hς����H�#��>���5�"f-��� �m-Z�dpL���3Q����7�}��՘���>Gky��������'!��q����[{?�O�=�Iw��+�x���H� ���W����{\����sZv���l��`�����pV��|�~���(���)\m�}���jm��i`Lv��r�D���vdE��y�(s�����\1�^����i��X<׍B�3wj�Il�w[�Z�]*f��H��y��8}.��f&���C�o�7R8�c6c\H,��ŠH����I�����Y��.K�tT@\#S����&X�<�tQHy��9Ά�?+>���jP��Χ��o�3%r7�B>*����t��pbe�)�X�b�S0���~�kVO��b�0���+���-��gfD�.2���\��E�2Ěԩ�snqq��x��1+ZE�ٲt��ND�)f���J��n�S��0?��>?�kb�8bZO�8羅���?���ܻ����u&�@�m_�7?�u�zꊑ�fYk�,av�
F�"�ke��������oO7z�ǾE��B�έ\����3L	�N�=��M`˚b��ʊj<�/����W��u_���9- ��D2�ͦ1v�x����E��:��Y#��]Bt!6
�(,v3����a�~CLDƵ��@F$��>�R�Y��,�`�A0���g�#�%ѥ���CI �O5�y�&�Y����.����P�v#�,���L��j�?/�6KO���B"d$F��~�%��n_��Sgn�$ ��l�=�!ƫl�S��"م�o�:g�٠i�	�.tn����&�S$��M$��Ɉ}��F�&挘0a�ұ�/���9 ��\�v\g_0�8�b)������E�h"X%��Hj�8�؜܃)��0�]X1�Y[ˮ��F���=lm�����r= R|�:_Jd���W{�gJ>��7Cr���,���I6�Y�!-����HBD&�- v��9}�L�q��%7��d1g.v6q�R3�{��n��*�?�޳ǲ,���<o��4UYY���ڍfDb�H$`�/�`��G�@i���D$qDΨ5~ؾ����\fV��/�7�h��Ϲ�FTvs���n!*2����s��{�m��0��ܵ�,�o4��JN]��;/�y�K�,�>��G���5y�{�"��a���c��#r�~VZk�G�yq����s�_ε�\fӅ��B�����s�ݛ�������O*��|�U��e9�8�X+�]_�nwU�Qӄ��9����e���_UB	$�(�b�5eA�5l"R�)^�e�"7$7��ؔ�L�����2tqNnV]�T�D�)��JLN�q�M�;ܸJ��Y�S�@c�tSk�Wq��V�8�$Kj���P�7WQl�h"K���yU%&(!�����������A��4�5�:���ؠ���d*��X�%��AqE'�Hm�9|�Q��K���}ii����\�_�i)���+°@yt���P 2Y���3O�^���9��T�l�,oay�2�)+�e��Ud�#Gȋzb�dR��j&�tn�4��2y����D����7�p��Ts2��r�7+�	Eg���\yV�b�Zݳ
�Ȱ-+?'>�ѿO���_X{��������ϹD��R�Ќ���ShJ�FN�m��DG�u��>v��.y+�L�+��:c�ӵ'f��K�R��Z"no�R˯"�/�q=���ٲ�%�r�_�8���Es
����d�$p����ZVzI"�rV�t�P���V�����a^�s'�ʗ�x��"M��HH41�)5�d6U���$���3��[q��V��2�*�f��8f&��؄2�l�_j�Eu���D�z�ͽ����=-;H����%��+�{�<\��LE��d�eŪ��8 ��E�`��tV�)�U\p��By�P3�Xd���QN>3a\Q�N��n9N!yw^�cYGʰė섚��/�2}���j�<�t���ܹ^�s��p��E�I�;���l��%��g��u<r�Q[�QMF
G�5�;�.�H!l�a�\�K��tZ� �����hص��D�4�y9kX��a��Uj�aq����i��L�����R���������l�)q��5���괳���ݧ^ÅK�~�̅4��C��%>�gA��@��"-���W��[��������X��\�<��������<���t��# ��~�j���UC�(%3�M]5���;��B&ʭC�Ue%�}%^!�V~峈Cˎ6���K sFX��;D�1h ��XΞz/T�����ƟC�o�*�pEקr�;�O	TDD��Xy���/4��V�2�8��n��������8�ս*���&׎?
<���W(F��yoB'���u~Ջe���h���Q��G���E����U�1�ܹ�
�^`n��������m
%[���wY9�q�����s��e�j���v�������4�\\�)x��"�Z�ε���B���Zu�����2A<�8��{�3��u�<��Q	"G��\�����;y��!��i\�\��t"Q�Bqh"�{D����h�+,��r+�Q̕�@��h���II&��ܗY��cްbRղټW��qf\�g���Țf��&ru-�����NX�M�ո��,�G�u(���Z-��3�T¸8�G��0BK�s͐䒞����� ��J\M�pn)����'ӽ���i�����hl�6�ޜ�I�|��H��#�B��psEo����a�~L�ص��ڱ�G���p�Ώ �
���_�)�>le�"-B,A� ���/���p��N�2,�&��������׳Bب��JN���M���_��:Q�<����!3}�#ɯ}��w3_o��P��{pB��y_w��1t��o�5�._K,�2Β@�M�Y*�k���X0C�	�n.�n�L��./]�gc����
�����$��KX[&Be��u�]����^��ֻ��\�/a��T�fn�:6o0�x_�/uR����zm8��d"wo���X-(�XxS4��ucno51�%_q9�&wY��-�@�NIy���z�%77�C[>i���qOzbB���U}ňq���j�Ћ��W��R�RY�_q���)G�.^G��?\N��qrn�'�5�h��ԽO�.g8hvE蔡�����
.�K�3��>��k���B��%��#�Ǳ���d��/g�0t>��O��R�c6z BG�.ϣD$�IS��)yࡆ���Mn�_�:H�*�-��*��W��e8��gD��BC�[�5��a����Ս+��,>bB��)��E_tG2�5��eew���B�_/����;/�6A\~�?=����(+�EG3�%v^*̼T+XJ
)7��Qc��F.���S+�S0���Š '���+����B+[
'F��O�:wgnY�lU�Y��u��>iY���/�����R	Lnq��g5W�`�P���8�ן��g��2�K�$+���,�٥���q�~A��Hy�����������|%�s��fd��c�O-.4����99"�b֚�D����eg��*��+ S��b=�2�m�ۘ��M51J�Z��2O��YUP�tsUQ�fa��g��m�׈��^�c��@����1�j��ԍ<�dd�����:zհ1Cp��BG��������޼���+ٳ�S�+yC^��W�X�9�8I�Eᙈ�X����$�B�_���f\�N�ȃ�-_����T_TZ2ޯ~��^臛_8�Oj*��k)Ă+��(ץ�����ೢn�+�n ���1?ϱ[ �ҸMy����E��塹�]$�@>^�-���_V����g]�zV CW�V���늵�ܮ�L]U��(�Fq��� &aT���'t��<�������
Wb��
�C~m��Vr�@/?c�X͵�n��dK�C`V�y{q�W��t���_�/�)�����g��5��������O��� �*_��������թ禐oX\c�3.�sj� ��r_֖�$Co`dK�)��GqY�b.�[�&�V��G�����9L��{2�_�t2R��.f���{�
\%ʆ�?OÃ�Q60����~�o��f�D5��f���j�^
��^��q�ڞ�Vj��>^4�Gy�^W�C�a���C��E���.�(���=|��2ғk�<�������\W_���K��7�������_4�?��7rUqe���b ������|���+�6i>�zd`�*�p)Hh�UeKC�J,�)��Tg���=���ב��~�5POF�c�~��+K�"��>��X�:O�F�c(_�+��[���F��NKs�Y��MIQ~T>���W�,TI��9fٍ5b���!.�2��e��&@j<=��ӈV2�"W���;p1u�:��)&�����)F��;UKJt����%-�x�ߵ\"��اf�ڡn[xc+�=���~.=���,�s�g��g$+�]����V�-��0
??�N�E"���s��|݈��lJ��b��Uwr.x)#f����pȊk����t9~���^��Z�h�<xv�)��{K�#�r������8Ĥ����G��@RK�(�Дˑ��v��̊nI&��/��^}��;��S/���ױ��ҵ��P�ܓe%R��k��.+?Bo����_$��ˌH�/��Ȋ�~�J��3]�C��7(
a3�p��*T|�ͅXdk'ZzP<�t�']��6��/p���6)��^�|��=QD�Xb�!Rw�̟�����di�|���J�qr��ųb�{#�.�帗I�y�Ng�`cպ�����w��C�;r
���Z��R)2WrD��iM04&-�NT���=!pe7<���S����Q_�x�U�H>?"ˋ��l�p�D��W>'�����yb�����{s��hP"�8_��5��Q�������{��z/�;o�y��J}�6�?vjc�?m�[�U-6ny�q�.b��Vp}$���ν'�{���(� ���t���%8^zŋ�_��p��Fhq�,Y�B�8�����f��2]~�J|J_]&�ؿSG<P*��"^;�K�����@r���:����Y���ֺ�����s7箬f�d���+�fG7k�-=Cn��>�i��י��R�����N��)�����)��'�H���<K�3�|vt��C��38��D����6M�"��^�Q�#�놆C<�!�N��E�x�5��C&0�R���-��+�s��ucˌSS�qa��3Nm�h��D2\�q��v���V�D��[|2�iRs���ٳ~\WK��+H���P���k�E>�6-)�R�;/�v�¸�6M�����0�͍�;O�3�umљX���eSg+?R��X\񈨙�/��>��>�3yA�Xx/�K��5X֒��������^�ݕY]]���V�����Z�ݠ�`;K�3G�0w}ο�Y>#��W�%8^zŋ��E���P��L�۪( ���!.�FTR����nR�/�	�Y�\�$���G.1�V����Ȯ	�������߿� ��2d�dW���e���6��|��JG�!��t�2��\	PQ�q�zR�l^y�������i�����sԽ�IhBͻ5	&����f�IT-�*1Z���`ȗn��|_E�&l��B��59'R��8㟫���'X�����nM9a�p�9��|C�m)ZD����S�~7-)���ҐPqfL^�ɔK��g�����}���h;ɪQ�� ͠�$O���QR��S�ΐ�x�s�穡�P�P�
G�@!���z.!�ex�����E2WÂʑ��������h^�<���w�-
ٱ�5��=ǳϾ��K8��dlE�v�xf�Z�8���C��ֹ��!�[D�
���)MDR�+����p="U��$���S~���K�]�&�˴&1�3��d�k�z=������3=0���띰�'���d"��}]^{�5'�H�����g:�^Y��YȋPV�%8^zŋ��,+���|Q|�|p3p�qE���NxV�ǜ�n@I�"a[�5�,\�U�U�f^����_��Ps���s}���)�^`����E���^��=�G�w�t�����bkAf��֖Ϻ�x_Z��b�A�mx����������m���$.;9�W�	�R�Sx��.x�,�2G�*t��2�o��;]_܇2ey��e�.p�66��o�<$R�����N��u�����?��w��Zݿ�e*�y���G�=��ACE˸[YQy�U���y�6��U-�I�B3�$ƥ��-���9<J��S�>��������,i�lY!�/��7ru��,2�i����r�.b��S�{�ZDʑ�wJ�=�p�5���l��iOC׵G�i�y;*�P9�I'�D<��1K=)��������bZ��u����E�]����j��H7dW���n�Us!���`�]M0uF��u�6~������d�����,�>����
Y�fp�1���Z'8�w8^k�!ڐ�?��bS^��W�Y�U����fb��>g�������X7'⠐���h*����@�����c��k(�]C�8^9.Ǚ��S,�گpÕ�����e�0�J*���uue�^��\ q�q�E�(�4[S,���2R��fY�������w�|��x����)«Ja�@����(���3/t�c�e�%�2��
f�$7��3�{a�$��@,�$JnS#�
����$�.n���v�����+��'i8q�4%[ދW�K���{[�K��!Zfk/c�L���<'� ݜ����ױ7�"�D2�V�Ⱦt/̗1�r��W��S&�p�|}'�9�&��(��Uڥ�/;O,��B�`]FN��Օ̤'.y+ԀZu(��b���Q�O�&L�G�ר6�Nٔ^ 9��*�c ��wL^�X\s��Yj eI\�~��3^@��[���C~a,Y J�{�Y�l��	����1�n��Wr��֣FA5V#�
[]��~�"��7�d��e�f&S�%��t6��g��d!����:n��z#�ǂ(z2�ug���n���_|�j~�0��﮳dA����a]/T�n�z�n ��@7��rpc��%���D�i�����I��Y~���s�u���?��:/���)Nb�#1�+
5\*���2(!�+�@\��Z���3^�[�n�<[��8W�W�eeYa�SK�C�'��c�e���ʬb�+ͮ ����;��;s5���D���+sRVb��q#�Vu�#K����X[�������+U稬4ðp�� ,�Q��!_��}c�ǣ8'^ӯ�ب5�'�R<m��Y�$��d��M�"�l�=)���ܸ�-Ob銍o�g��ԛR6�<��f�Ư���'D��,V��<aX(^��c�5��(U���i5�\�W$�q�"�j�̀y�)�j��s�8k\ѽM�t�J+�a�J�kR�d�l%���:��Ê61
����B��cFC#e�Őn}��
%�X�"�r��qr���e�rL�s���yS��< ��ڍ��� �
w</���.��*_�{|:.��(K�z���x[�v��9�D���]N��K_�Թ�Etk[Ǘ,�*'z<���v�I$K������Жi�Bf�&订k�aF]��T7�����Z���XYaf\��ŕ�?ʊ�,l�d'd,��^�K�p{s�o��]���kg��\W�<t[���n��߹�%�.�E�_tD�1��]B�v�6�`9�°������%/�}ӐK�b�xs��ϣvs'<6��%�e�W�Εhn���D�>F��h��(�]�Gm�x�8��N
c��-�ԋ��I5��B/d�i�2�ϊg��lZn���آ�ڑ 6@ɿ���nQ�}tLX��kT�ݡ�;R_�w��!dU�UR�\������b4��b3c�ʭ���H�8Ş9����^�+)ݟ���sF�9M�=m����ȻU�S�FsX�4��<+�I��f���zE����P΅4*T���!s=�kD�c�c��a�WIڃ��"���:�G����W&��w����po��C:��8��#刞�R�5�(c�66��z�E_�<��V�o��:�n��\k�5w�(��������rvr����z:���h2��;��������++]�S�!r	�!�y�}־���Ƃ� -���^�E/���ԕQF\��2ˌ�M�����o�l6e��LAɅ7������*��'�=��d<�Q�R��K��ƅ�zf�?|l�,���9~	��6/d��e�z��r��u��]��]龴!��\��>�5MJ~�/�OP$U���_�z�h�졉��{�+���;Wc&t.0S|�,���<��UY�͇�X�ls���%&Fbo�>�I?^�K�*u��W��,+��+�|rE_�AFT���>jk��e⒢1.r�`�;)i��|(��\�`-Ӄ��7Z,.� B�p�ul���u%����m�rIФ`�[]���n�I�j�sS�L �����R�ݍH���Ui�:i��Lr�P�k�
5q	Me�	^?pno�l�R�<��
{q4.h"3&#�SU�|2��T����t�b�bl@C��Ҹ*�˹>�k�"�	�q�1�>�Y�͎��a �F���a�{h<��r6�J6�,n�s>�"�T�ry>���>�H����(^�ʚv�J��?>���}�V�}Q�Vdp�S���j��ޖ�~�5鬭Jg�+M(��ť<{�LءmooO���o�o*`���g������.��S�l)CIS�p����ρ�[�\��$1�@CHq.Ӯa�4�M�C�E�2XaQ��ReUTF��ğ�zU}����1l�>b{Al�a���5�!6��(�e�`����]#��Ì@��_RR��0��=e�!��3$�����,�m��J�$�=�Zޛ�c��]-'�ڔo�h��M�g=*�N�Q|_�a|�4�+W�Sge�=����<y��푒�R]rT��O��^�r�.]�>G�+{d�C)�r�ݮ�f��}X�P�D9}�5��q�.�ހ�f�mL�[V�A�q�;�m�[��C�Ey����1B�V�J1Wi����塙���"N�X"�Qm�YSs��]��Z�/�bU�+��5��S���Z|]�Y�RI��E�i��1ύ�jV�`�eY�ɕ=I�J�4�.A|���L�<y�ٹދ��e�ρ	��U�D:5(/U���7�e1J<K���1�I�1>�p���S( j(��nG6��2���ڐ�|('�c��3	[���ޖJ�*�ͮD���yrt!?�g����u��u�AQ������&7Y�2�nC�6�rc�u����G?��%2��ǲ��%-�����|�w������]�X�x�+7o��Ζ���we}sC~�����h��ƍ����k��|R�����rqv��ւ��0�<*vXE�����]����>O�7z�ϼ��p(ۅ%�5�MI���e��p���{O=z����+:�|����'G���ɀ.��}����n`1%�"��e��}��5g�\�\d��W1C�sn
%ue+��Al<��+x�b����S��ʲ�P�z]�T�8�h��=�kZVm�[M���OSC?�(%݋c�6_�(p/�2w��&����Џ^�M� �<�9����%?��K��~������״M�[&��[�����1�AAPi,X�q�J]��k�IK>VK�+�.9��f~43��@�G�U�k��Z<iJ���R�]{�k�+YS��&��V��k��I9(��X��K�Ӱ�[O��h�71pq��&]eο���:�03�@�F�Vr �L����OS���t↢�$g�K,���j"�Q�G�d;���8��l��υ�)T�\��2�>a�M�Fk��l��ʍ[��]]U�R�����HNN�8Z�r��]Y__WaO�,�{��ɧ���;T��6�9���C �Ln�mʫ7o@	tegsUv���?x(�d*�'�1kZW啭���TTx��O����\M<(�j(��t�]y�ko�����#q}�S��ݐ�FC���Kmm]�I<��^�B��vd��ʫ����#9�����@�Gc	+x&5y坷䷾�u�?�.���P.��Z������o���ȏ~�C�7k���:<;����w_��7o��X��_�{>�i{{[��[����� ȸ�̌���Jx�^�b����ʕk��;0��!AYӽ��QF�l�U� ��W�U/�Q�VB����d	���#"S�A!���bIx�nC&����ZNgSib����Ǡ4颌#,�y�ID"Y%�LD�k��v9��g�b�O����#�����[/d�p��
Q�m/�������h�(�g@�vK��ܻU3H�6��GUmc>j|Z�fd3u$��>�T��Z�1�j�(ߨx��F蒈�f���KV��9�
�ʧ�A�P�k�QJH$�mA`��x>�Z�S�&�4p=��C<�fő��'�hUהI���U�Y2�4�@p�V�liFe��@��=H�6}s1��i�<����R�u:���"մ)aZ�hB��r�F��s�|,��D:�c2���볜N碝԰Vhpq\�&�%��Mm��Y�	t,� Q}�ޒ*��I��E�P珮?�o���L�g��T��:PW�a<��9L �O%�̤���؀�!���dxN>�Z=���u�b���8#���ٱ$��ͪ켱+�- �j�����#y��C(�T��7��s�J*�].������1�斴�nb=�ݹ*�ɬ"�Y_��ϭ&�������y˵~tBeUdcuM��J[v��%��jw�һ<���mElT"�[��|9w��T��)�~�1涭)���~�;��g�@1_�͝U���w׶��ekkM��[�J�����H��-�dc�om��;�#G����ҩ q��۩�&��^k�?���D���oo��,�Az)��0�щ�w��-yp�X�FK��r��V1�:����.o}�m���������w�����R�ua�U�������zC��[8��?�H��;_�^�����敼�֛���O4G�ϻ�ym(��t���K@��9͆ƚ27|���ޓJ%�:�0�d�iBS?�x��{0�Υ�;UD��k)Rj�Tˑ` |��'��.P�[7a��c�M���%8^z�;K�`K�r�EG�-+�(uG+I8ݝP��Q�LUT[3Y�*�뫒M�R��f��t�=Y�.7X��H
�N��.n��,E�yV� ��0
Si��9ΗͪP��
�80�fK��k��B|�V>Y��肷v	%�V^����1.Ԝ�=U%[�E�q B�D��"W/$K$�P� �1�5�RoU�K�P=���c�����X.�	���!�.��ͪ�k��&6UKb�����H�a$)K?�[0R:��:�;!X+�+B��h��1M�n�:��J]ƃ�a�,0cV��ҁ�H�<2���B�H>9�Z߁$m��f�٪v��p.= ��nu�$mo�8e�$�,�Hr�X��4e��M���P63\�,p�_E��*[�P^����[Zbrѻ�G�I��[���l��r�z������'��ߗg���<�a�ŲVS�	 Ԛ���r�����U�m~H���>��!��L6��e�܄����%>�및9�lv���
ƌ�7ץ]��@�Ai���hu�Zͤ�cc��je��ݐ��X���ěIp�խ}�M O�emwCN����ߖE�"qcK�n�.��9��|(�d$++X�"�P�w�
���!��9_x�j��ػ���>��T����kkk:w����{������Qqp�����������U= j܅��Z��j�ޕ7ߺ#���i v4����c��`P~�[�ʏ��oe1�ɷ�y[>��3<m]q�	O�"d�x4��ߖ�c�g�[]���ۙl�r����7�����ō��zT E��`P�
c��Y�!滽�%��@�c|��"�^k��9��7��{���٣�X����[�M��s>{�	cUE��sW�L4]8�ꁉ'����ŵF��|�����%}xO.��O��e2�{UWV�s�뀙�4��z���*|M�Ê��K�x�8��yA�p3RmU����$�q��-�"0lC� �d�9,�6 � V�l�Q��r��Jl�[�E�¹����t�� �z̏�5d�` cn@(A�|��QP�s(�:�L{�N}:W4�g��"����	��Z�s�x>�IއbɈ�p� (8s�ĖM{��Υ���!cq:-w��'�T�P��7^������ �EK%J���{��&PÖ�#��g�'�)�ܿ�˿�ӃCEZ��+�0�3�8_5�5՝պ�zcKQ��!�8/����SY�9��
;��-&��.!�b%7a ���b�..��:�a_��h��Դ�9Kc=T�w
�;�B���5Ĳ?��-�g��&=(����Aw�J�2�Iʇ�E�K�����lDMYi��~���K3�jE�.���B�uT���?��:==�d,��/��p�ލ��G�U�u�Hk@�T O�>���c�܀ �����.���JK��|�>�evٗ�?�-\s�kocC^{�-<���9�Bm�%�p�u(��;��i��&��(�%�nSVW��ހ2l�`���޺4�~j�t�:�������\֥wܗ��d&sr C1�5�{�O`X<����<W�x�Y�3�����������gR��8�`�I�e�H���鹬�n�����\�&5��g�ƾ~���)Ce�X��+� 	�C��A�z2<'����"g�?����ɡz�TJ0�Ր;�+2:I1�U��4v�:�`�>�N{Ͻ�{�л� E2��R�=Zuv���ƿ��)���d O�N0O5I k.��G��$i�hE�=8���2�=N�C?�3��^���@��o�N�f�/���\Qӣ���qn5�Lx�'��YFy:dK����F����h��ƹ��C���O?�8W�:� |����h5��S(elxn&s�������p$Y�[`sf������;�L���P��V����c�P��~���W�:[����k����f-��U9>���?���*x-!����bk��,P>�] �j�.g&��{�KI@N�UY�AحWd�1Oe֛A�@�,�ڱaa)7��@�M��`E��h���b ݍ-�U(ts%��g��c�R1C�o�R��Wd�]P���>�r\��{7��m�=/cmDg�;�)��Y
����s���H�WW�h躚,Z�܊�Z�����Ŵ֔[T�D�krĊȓ3ل���F����E �����r9oVp��o���	xzHk�k��S�BH�Ԡ|���B>��6P[��ᲳӒ`h�Ay�8����-`�L%l�%#¨c|�Sh���!�N L+��ii�ɍ��,F�>ƅg<I���
х��Ɔ
���ܹ�8g����p�`�y�V��{��m�|���Ԕ1@��H��vp�cy������L�ѥ��n���5e�w�������b:��xfa��zck�"7�x�<�A���֪zM�<���"�>�1�ޒ��59��謯Ȥے6�٭����L.SY�yC�#(��u�+��ڛ� �9~xO�b}���𳻳�h��7ߖ|>S��^��Po
��nhЍ��򳟽���K]��Vi3+�y��w��,�����)��#Y�XuT�������l�ۙ����f	3�	d�%r���IVcJ���7�02����j|����P���T�������zahh�1��<�KI�'��c������[�,u3ɯ�4<�9�֯>} �ېjsKr����O~�Xz0g�D>��u�7��p�1��O�S��D�7��/`,�X�ST�j��֪�"���p�J#��Z�֔���(j�NR�\�5���4�{g�Z�::Q�r�:?=S ӆ�j(asQS/3�Y��^
��R��o:�V�Re�	_�@t�%A��WZiF��âۀ0Y�><?���E�߭�u��Dbx�b�r���M�Mcـ�&��h$�؄0�������&�¢d��Io��!�@2�߆q�
c!�d8�b�a]�.$�P�|ݶ&��P���*��X�9,���ܖI��F� �4,�z��݁5�TA�Z5��M�]�N]��ΪT;���<Pi���ͪBߥ!�%��G3Ғ+ k���"H�q�!�k��ly�������P��:�.=,�6�B�~�_�|��^o!&Y߂��� Ɠ|A�ޖ�EO�Q*7wEj+��d}
���{]��TN�j�\��\ج��� 93���ږx�
$�E{QJ�I�CF,�@��o�Bs���y����;�Z8ce�#M_���8R�9�;�pi�x��P���������=��t>k��Y������DP"��ޗ��'���#nE��<S�J��ve�����`f8�%��&ƶ��V����?�u��ܺ�+��H���w����g�1�ɚV����ɓ��|%����zK9��Νפ���
�K,��5}�s����MyL&�$S/��Hnk��M�ݤ��P4X��Uh`�4sJE��f�ψ���������<|��T��D���/aTb5`tU��N�d{�	_�0n�E`�W�҆��}�P�g�%��3:m���~QE�{�`��p�Q=�_H�]W��Z�d��K�[�!����S���s���]��wHC�(����y�&�s����t���lMV�xև�����^�!�;�Ĺ2��4�l����*-S�L���ǵj��oB������ʞf�Jr�3ǁ沌��J����jx�����B\���CH�Nz������l�u(Cck��Kp��7,�������� �2i�X��tN֌���*-qwY~\�L�� �u H,z�A)oX&3�2��չ@�K��y����9c�ЁL�Z���FA�
avA��f ���e�4��dП�CX��t���p[(^(9l��E*u ���H�t2� �}�
���iA!�'�LH'���(2%C�݉��}&
!rh�~ʙ̜�㿕��HJ���RĂ��qt�c�b�q,Ӳ��Tp�@�㹎���X@ ���P$@�HX?��w܏��:d>����-X�PT۫2�(�JGn|â�{kJ�5¹I�P�㹲����[oHB6� 
'9j*)!*r
������f ��P; ���o��o�a{);[��n��>��B>n0a�p{_�?����]ZV<�"8�����Ɍ]&�yf *��}�{�t���}�{��dx��0�N�5V����)��{����/��â��6W��M74?��㞬T1ߣKa�\�5�X���!w�"'�����̬��P�H�r����d�N`@�e�-���zN��9��,#�������D��ʮ"9���ϱ����U-O`$l`�I��D��M#1REJ���mP���I�(�:��rCq�2!�b���?�(}C�3Ě��nlɎ ��h �x�	�k����_a\�!|vp�F�Hbȉ@��1F�����g�{]���ʖl��M�c�r�W� �jveߋeFpL�.���3�Y�1Y@<� ��{�AMv�D�_�Y�j~�q��)J�44ʭ�܇���}�|i��$+o�����s���\f��*��n��\�����5�\-d��J�����lXP�k+�Z� ��3A\���:^z�+�g�?�y��KZ7f�	�a�q�hm_��(7c�sY�B{v ������
!톰��*t[S7�|����Kd�ڕwn�",�&%$Pha#�2�do{hd��K���8��ضMI[mI*X�L��Q�Nu�E�(�n��B2�'�$�]iפ���a�kV��f)PA=m5��}�p!BB�jE-�6�C^�f�M�M�ƍ�4����@1���#1n2*
�6��[�K��gf]C����������&���wߕ��Rvoߒg���3���M�r�k��������?PT: ��"������;��������d<��
s�C��Wߖ�7��pp&YE��Is5���\�7�[���\B><8�$�g�Ϊt�UX�k��~K>��ϵ+�{��I��綻-k�+ʒ4�b۹eq�����ּV��70?�{hU����L爙�DNEK�藊���S�����v������V��g{kC�0����^`-��`��ｭuY��o3VʵFW���<�\�u�����|���H9;�"	5ƹҭ�Y�fBW�+0����ˤןj�z��[Ե�zyvr�Huփ�r2T45��*My�옅EZ.������C�U��RV?{�\��-U�DUMlS�/O�@�@�������X�-(�:���*jͲ�{��ӭڀ�I*D](�F<�j����Z��'�9%�3e� �U�ʝH	�'�UP�4PÐ1�v��[�`6� �B5�2w(�V�l������o�u�'Joɺ�f[������4�9�3<K�=sl�X_���Z�h�s�!bo�H�m������a��0驳���\W�)�Sm�s-*;|�oH#��O��;w�ʽ{+/�6��������'����FC� ��M{&Z0��}�����Mc��ܸ�+��Q��=�R�_�#
`OV_9e���"Z��B�wdM.�	Sl>O�@Tj���&�0F�:���� ��c\���B�o�hk.(��M��w�#�~�C��H��We�6؝W^�w�{C����0�6z�&�`��@[[r��-��Bx5!Їf��A�om�J}o_�3%3ov*rq�1��!$����n�)?�H�%�VU�!g�)��My}[��/�AW��p�%N�
P�;_[��?�g��?�;�^���2v��o�`��䬥�d��0k-���P��z�?|�l_ܠ�d�;����ʿ�˝7^����0>\&5^{SnC93;��[�� ���-9<<�ݝ������k���]鞜�i0W�Ԁ�g����VC�@)��O$M��Z�C9c2���qkϟ�>���4�0�y=���R���7���!��z4�H���r�?7F�u��t[�ߨC�Fu-5��Ø�^nT׃ջ�}�.疆!����c�q(���L���&��\(�F.�ǚ#��@�{2�غ���40<���Oe����d����8c��Y���#B# ���@�#(�Z�lF2�aoLd8��y�UU�I~�)n�F	��\�Df:�F�&3��������C<R�C1%Zu<�����Kc���.��rc�2�S����m���2�Y�DŖ`��<$:���]@Q�jʨ�kW�t�V���z�j�ٸ�Ge9R�<!ဟ�<����	MƑM�d^��G�y�:X�L��+}�O�ҹX;)6�|v�%�ؑ�1�%aq�uݰ�zU(RX$=�V2�4�!,>���zc]va�_<}�׶�I��ŚY&1�w �5�'DK&<#���H̽�=����sݨ���d�b~�kf���Ho3���yN�?=_��{#sa#��N|�%;^zŋEik���PQǳ'O����*����Z��
5��S[Uݬ,S�c7L�.�W_�����S�����I�v����i��2��¬��oܑ_��WRR�{�,Bl����[�z���g=Hy�&���L�ro����]y�$�y ˲��)��@�~���z���i�oɃɑ
M&�L�UiuW������_�� TI.`�_V�FcGFY_����+���&>��yS~���R��ق�]o�q��E�p��r|p��Ϟ��J�ڎU��jj�|�%S)s�}�䱴:]�����G���s�9�~r.'@J}(�*�׾���q|��l�Ve~r�4wd
`H��> Od�ƾ��D!O�����Ƽr�������˺�\Ά`@�] �l�m��ۻ7��O�{J}�l�ߑ�����8�t�P�3"$&iA�������_A�~�@rs9}p�(�J���s�^�Ž�r�]e|&H�ۍB�{�cj<�M��r"�/
8�S�������އR��.�x���ǵI�G(�J� �=z�5��7���y�al+8���C9�5�^�)��:�^
�g?����74�L��FѢB���XEe��1����T���J���r$�������j��L���sf���{��t�4�k��\Q�/DlK�/����xW)Q�J���s���@�^���J�Ť�5�c�=#��V�l���9Rv1&#a*��f���%��j��=�:0��Hgg��'������n�p%�'Y���R�; vf�gs��ikX#y�1�K����ZK�޺bɟ�}[w���`�K��@f�+ՂB�y"�k���,w#ҷ�M�/��ö���F�rd1�"?���h�Q��q���~�����/��	Ppvv�I]��� �����"c8��/���B�D�j(
��ĭXf�h���K���џ�Q��l�eogW����]�b�Mc�a�^������|����������2NeлT7�ڝ۲v�L.�Z�q|~f4~l7e~��-�������w���{�1jui����5�'G�3�C��i3��IM��;����b���-�<=���-!oBq��ٖ��@D�ByJ�����k���=���/��g��H�Bn�vG�=Q��S��րth�6���QF�q�3��?*�Џ�cU(���U��?�wr��=�Dۦ����c�Z^u��|���*퓟�/C�у���Cy��M�k��:yj��X�6����)�L�ڐ�)�`s����zR�\��U�اm�H�&y����顬���$���@v�z�\>��	h,G@ߏ�G�H9�%�(��b��z�G�ޗ5&��n��J��9�γYX$X�su�>�j��qYnD��9W4����B��,+ʡP����P��1�%�֞��]*���d���.����M%���'+�o棾D��*8Ǧ
��*�v"U�I��>�V��v��[��47Eɚr�<����Z�%A�$4��lc�;��\Ÿn5��tm�j(%�j�Z���$�g��)y�Xx�/�Qc�c2v�x��iH�]5S ����0R�/Lr�ђ��Z����Y�hs��dR��5�U��x��9����6�ky����J���KM=B'��I�#]'�M��6����ElMYBSp\W�!0:S�9��AC0���#�$7"1�;�Y��T*sk%�� �?�k��U�H����"!�{l��z�d(,�\��3�9cwE��"UCT������X8��=��O��p�_^@�u�Q�`ٴ^D]5�:kaܲD��@E�2>�H¢�X��?���G@�M%� �+���؏>��Jvܓ��u��������'�~,��z?��ξ�6�dr"����?�XN���5I��2崆���3�ֺXOT	29h�v��g�Pw6ߐ�������@�.�����w�&g��������'?��|��ϕo����}S���'�7oȓ�Gr�;��h��K��ew�����Mа�O�W��܇~����⯿/w���ƜB0��3l��k�)�<���d@L�PbU��\�Tٺ�B�B8Aa����c�B��si���e���H|v$k�P�˱4�@7���s�*�iĨ�T���S�f���w��=9�/�` �h,�2�=�=�w|�P�� ���l@�N3Y��68<���X�XG4����"��nG|;:M0�����O��3��4�� Ѩ{n:SNb�;��RcV�0g�B��b��r�g�qɀ��ĺ��f$kɭ_,y��c��<Uv1b>D١�v����5+%�k�Wg�!C1�M3$G�� �0���B��"B���Y�
��@P�Oa %in?IV��#�[�=l��G�V������r^�I���*�;֗rh�SP,{`o,F4,0�ܲ���5;� ����,�H�%��^[��s]�m1�zғ���Jx�sB�0���8jm�b1Ř�bͳUo�$�=R�f�\ۊ���{�Ơs�f��k�{�%�|X�p܉����Q��5�6�B?Of��C�
��>�1C��GJ�A�ͳ�s�9"}��En����L5�Li�6�ZUI��Q�@��Թ#2C���7w��/����3�A9��e'�V��m�<	�A�Q�Mj����F�[�r�衢�H�bby����_��\������=,�XKd��$*����L���H(�\Lz��)����P���' H�2���dP�IGkp)��:�&o4����"$!H�mpY�K0�g��%l����"C�={z$�ˑL�U<,�����_Ih��s2�"��`Nf�ҕ��b��f����OY��1Q�0�����'|���?��m����ӏ�:��0�Y�=��(�>�9P��{�ͥ��U����}I؁����_h&tDD9@i`�O��f@�@����Dl��z)O1AB�y(�32o" 6�{���Ls<�h*0ZokG�$�4����@bf��t&�l5�ڐ^���\���9��@�꠪n�(t|��Z���������P�2�Qqг@�>\�7�7_��-�[f�7�AX5��Y蚼��x5��d�����c&p1�
�wj��a�	熜��\ϳɬp#��L����4,�{�統�-���Қ,��R�Ҡ�[]ښf8�5�1�Ps0�f�K%$�.2׈=-ܕD�i2Q@6hN%ݱA5��s*��eI��ͬ�n�i��BaY��;��JT�IQU][�X昻1�0��4��H\�/W~�U	Cz�&�+��J>#f���>�?k�3O������)M�hj�%���w����0���!)`� <����2�SvA���S�:c�{�믻�(��NՀPT-�=��Ϫ��f��5ø��KkHv���al7��TK)�eq_�i^�T	c*U� [0�B������#�d�W���~�A��&r%ӭD���ZD�Kd��Z��U�v�Qw`k}JWRE\h�)�3[�1�����S]@�@�<}~�M����ƶZ��'G�rtz$ǽ�f�VH9��[�x�{
���:�8�_��X�f��>�ാ����Ca���@IR�F�#l�秧2�f"9������#i�Y��j���Ǉ����c�7���!�Cl��ؗ��9����O>պa�U=���E�jR�̺�0q���|�>х�V�t%s#��c�ި?�����T�L0���[#�	�	J�	� Z(�O#<�f��ҟEl0�� {���?�VJ#���D*���]����Y�e"[�`U�ZWŚA�N8f���N�Y`�����^�_P�J �� )��ؙ�1��jW#��H�m ���U)8�n9ESr'�|H���Y�Dk�w��%�Z;�8��ZK&���l���<��:������dx|	(M)�ϸbܩK{}Ud<�d:Ѧ�i7%ߵ=s��1��ず����uq�ͭ�]<��wI�/�(Bȯt�@�-9>�bS�`��@G	Z���������CE3�T�����6�ʧX}�*P�׻�>�o~��՘H�6*<���03�xN:W��\K�d�Z��Z/�ؚ��8��%՝cG-7b��f�-ڃ�ߋ��fnr�^�T�NMD�4�S\��_6��������J�ʮTZ�#\s1���p�4���NǓb���e6�����V}�\nIyl"B$��9��ia䭮�h=��A�\�e^�Rq.�X�bI�ψH��k��ܺuK�~�ӟ����*�rt��|��/���+^zq��^M5dd}o�@tq`�ҭǸ�'���\�3"&���j�h�;�x-�H��L.ԅ��C�V%�1��9������>��%��M[��`�P*1���)��+,IB[DRoQ@�]��?ɠ�޲mu��"n� PgP4�X^�����%�ό��M�#5��Bـ`x&�LF�������FL~ �n�65�c��zg�r(- ����
/���+�~�ڳغ75+m��mb%��tF�	�$�̵��{D��1��LA=g�:�5��I�ܸ�)$C�}�)P�۵��S!�l@�]�=�O�Φ
�PƘ�	�C��pC�TP�(��!4I+��xx�<7˲rJ,����R��-^MF1�;��c=�FJK#�.����+\}����5(��!/�^je����?��wv��Z�Z$X�Z��D�Ԙf$��7��Cy��1�m�/|A��8"Y�ݑ���2e�X9?L*LE�&�؄J��we��g�;�)鲖�zC��M�S�r{�L㝪�*U�.�w9����>��%B���Z3��*�T�:*ۑ�5z``�(�F�!�ͺ�)]�>������}OϏ�E%�f5I+��Wi�(8������bͭ�־p�]�B��0W�*bݓ���4���C#y���Xg��Q�GD�|6V�L!TS�~����q�al/�PɭoV��bZ�Ey�IFZ���%OU�j1D��4U��X�Ɛ%(��{7=�c��Jv2�*��3`Y���h��^����**���*��iwdkg[���l�*_���<�lp�<���K~��7�(��FJ���?�X�h�[g^&.1�B&�c���"�ᅒ�@\��X{�F�B<S:�jLE�J���imt4�[�031��B���h��h���1�g�.*1�Dp�]��\�p!�?�rj�m��(��\���}f���а�7[[@އ�̘TJ�1jZ�ӑƯ�P���cĦZi�F��i-]^ix���퓮�aY�p��@�$���ӕ,9C����7q��J��{�!EJ�Hi\�����!9�6���ڴ=H�[Hg��=Mm�0a6w�F�J�Ad�n{��z�T"�s���t����fS6�KB���B��R:նt�����K�ʤ�,�8$�V����^O�e���샨F�(�֪4�k2�8��G5)�G����s�h/�g???��1���կ�s��w�nH4;���{ku�	O�Q�h0�R\C��򶦧s3�JgjO�;�,�:�I��+�"�`�\�<��ɩ*��u��ݓ(�/// ���ﺎM�m���;�����HP�F�Ŧ.�D���e^Pz�~O��~U�9C�h�]Ơ+U-
\�-��"V���.X(5��N�y=�ᥬTa�y��O���T�;����Pb��:ka�\�Ü�`Y�ݱ����3^W��lFJY�ĸ��)�VC��1��k.�����D#�-����vG�4	<3��5�f�l�� �TSR/�K��}�7e.�[?f��1�j�+ʦ��U�65�5��#�,�1� �ʌ�k��s&�e׭��m����InMU�]�\l����vңg�H*T�:#���/��%C�.L�W\����Bf��nn1���g҅R���+0VTg��a���
"1��Jf����f�+�� �f�X)9�a�'�h�nK��e�ز99>��G������ɒ�|�q�̘t%�T�A�!�:��`�Senq2u�J�/��h�@�L�A����P�&6J��"���s]]���5���%��Jg�HZ��-Vu��l7�g���0Q�?�������eHQ�m"UC �7�~��MΥY�4����\V`$������G��&��F��	!,3�U��2 ���T��ZQa��,�݁�k�I
���Uk�T}�U�z�-5�/��?7���L�I績�<�d�Zzfmϸ�6֤���̒�(tFx>$9 �/��֒��c;D�w���c�K����.��,?N1�pm��Τ����:�0�ų�:!�җ��C�v���P���?��f�g秎���eq�cK�#D/���h�b������p.��a� �Ř�fjSs3������V�y'�]�(dG��ٹ�'�_�zFk�H��i�0�O��J��������I*��ԍ�N̝��#4�0��dy?3�Ӱ�	��q sY|?�<5�N����+u.۰V׸�s3��C�N��?t�Zl�a���Z,c�{����"֒����Ȓ4P�(��	��z"]ЬN��ݘIy!�Ɩf�O���9��k�%E�Ōa6h�(Gs��ҙR,#��y�+��lp@z� @�	�����3��Y�f�F��X����J�4�Nȇݴ�pq�李����/>���ݸ��V������0\�2�pï��L,13>u~4��{�����R������!�u�H�tB"n�V�����%K��SY��������b�����7�яΦ�澣;U;�P�du{G��ZU��Y2�0γ�ؔ����%�W׍���X=�X�Z��w� Xx�H7z��
*R�*���4���H�$H�%/&v+r�����{@�Eu)s��ihy���M��(��ؘK�C�Lf�Ғ�^���<�ݻ���G?���j2�;!�:�jR2 �y_拱6H��rS��@�A\�K��S���%�%3c�.U*4�dw��	����t�0\xϤ�d�PBWq�~��`�߄����RI0?�!WR��f]�"ʹ�$�W��b��c�s��_i4O�MI��j9χ����?;;Q�&ۡ��]��T�FÉ*�I2���3���mx�7�pƠava�g�Y������V�JM�u�ɤCb��ۀ�?}�8��sCET�l�׈7���3���B�㙪@�٭wq!+{V��d66&	1�r$�(�W��fW�κ��T�k�s5p�+����q%�D��Wf7G��PZC��֪�lt�g�N?LS�
��h�������i����+�%�a_.�J�:g�fm��'.t��(�/�� �̬3��EbD��S�w�W0W\��֋���3����zZf1��-خ��!�L;AեC��{uN����r
�co��iA����E��MR����pl��ĵF���O`Б]rϤQ�����7r��>)_4��4�[���@�q��a�p�Sf]C܌ss�{�[�iL�|�����3����0�Fj!'��י�r|p&��>�P���P��L	�2L�l7��0��`<�\�e?��re��p��/w����~���֛J���z�Uc��i#�L��X��+��&�r$.x�c�u��s$n`&cN�4�lJ&fY�fU����B�,IM�*b!�ӄ`
4�U�@D�%O&c���g��X���vX?Jwz��=�+r'B`�<��$Bo�[�;9R�;�:�0���Ko�IH�%�0�Ɨdi�sA����Z��7��//�䈙�l���LIV���ԝMW�j3v�՘��!r��d8�M�P���P���;Ӓ�`��1k��M��@�{a K��"$Ȁ�����N�^HּIP��\�!d����eY��'OKĄ�d�udB�c��hГ>*�^^�<r�.��ԘWP'�݃�?Υ� ��$��]�����K(�<+�e�J#\���ω�f,r�+u1����*	�p�]�`�kx:`��T��x�P�Tݔ�C���h�9o�-	-��-V`6�����u����b=1Q8�4x�7GPtշP�XS>OR�:��~gKN��wZ2����+��6� �M���(������4E�$I`��pك��P�g̾'b���=�U�$� cS�^���S�[V��t�>�H�e��̀�5]2�~=�nA�`,�L
�51_0"����(ǤaL[Xo���D�/�`x�3�_f��
ńL����+1̫F�f�Z&���<jT�x#E�D�FbF�d4������ޛ��vVU�su{�ݞ�ܾ%�$� !1$>���Z* <�����+_a��S�*;�$6� ��ZRjB�(���雛��{���ս9���������{W~�wr��gﵾ��َ9�PS�����.����n�h��p�8J�����^'��eY��U�(�U�Љ�`���9�}�l�9�6����tՙi����Ō�+��|�(����	�L�$�unC�G�F\4��{�;�eC�D��Y`5@F�]�����a!8Ҭe�N����SuH��@"�}�1#�U��>���mC�#�pQ&��}x���lmhv�JX�B�A��>ϔ�	��Ad8,˟MI��)������,/���wc%V�Gɂǁd�3 �3���D�@�nl�#G3F��񹚊���	��y���,Ԙ�DU�R׀������eM�{�?m߈�]��#�aە��Y�l+���	�V�1�<�����S��U�>��O�%�@���3=�m=�p���C �{�q�H��(�55��?(EB�P��e�xCuTb�ߣD�~'Z !SF_��q`Y=��P�7,���;�-]����aD�wa����l$�
�O�e���Ն;4��2}��2@x@~�y������F8jB ��(����q$�fk�"!�]�`�Y҄�C��f� �2�Ab-�K3�/n�V�9+�"��ޣ�?�$5R� �ip���K'��]���s����Q[����
�+��X�<��R���O��R���螝��.� �[O 0
����(�_���ϺO�.<� �Nc�����4��f�J�e�u�4 ibf�Q-���`"uO��6�pA��"�~#������rWW��v�3�q&�!#���k��{��;��h]� ���a�
N�Ơ+���P����7�K���r���:�]"�)����=c�Oy< �}�Qs�q�6`;2D%_���x��+�U�����švC�N����:˾L��������Tcf�|�h ����̈s�ۀY�jEc}X(v�@���eB���X���:����v����8L�C��X�F���>�	����Ô)i6��PgIm�F�����,q�`���X�cd7-����:Y&�Z�>%J��b�c
�Xɟ�P����D�K��_e����Z�y��ٻ�d��ӯSu<c?�N�c�E���|i@��؅��.��L�Tע7K�}.�77��s3�0
�G����>��D/}�N�*T�$���2eI�5�=D�0tmݱM1��L!�3�_
}*zYɘ�rJ3�����֜�$���p\�A k��LD�j�n�h�u�3�����&�=ʒD�D��ḠL`p�c="���I�Y����\��A��[�l��f��@O�f5T������yX7}]M\����e#Jぺ�85����s/�H�-�����C��1b_�g�l8�r��Я4-m�Vw��˫GMj&|n}�pa��W�SW�c$ñ�	u� '�^3z��'��nu��]Gi�ˮ�'������5���R�K��N6k�{�e����t�<�&׸G��R,J��O7w�������S����24��>���g�����}�XekC-H��h�g�ғ�&����lo�L7��a�=�\�M��������ߝ����ox�|��;�=D�K�����r��Q����dʄ#j�NP��+^n���� �($T[kt�])t��o#r�iE�i�z\t�Ɠ�L#`_k�pa��0���xta��	S� �C1�T�E-����})G1�"�Y��wD1�e��$(�~$�����Hd�q����7p�Y��I���c�l����p�.���	;�Bǌ�	v(�!�ѯ�]N����ܪ�1 z�&jR�x��mY]Yԧ����6�txE�\���8�%d\��!+f����Jp���@$[8.��!!������2��P4P!
��	dC���9�Q2D�W?7�i�˦1�5��Q���`�K��B'3���:���2E���Jj0�qZpf-�%?dj�CU��D�	Dm���h�^7J�$�/��,HI��q�1N����ʱ��9.Hb d-���|8g�ͬ��VY0�_�(Z�3S4j���oE�es�z�x(���Qq��P�9�H�������&�	c*�)��@ ���:`d���=�'Gй&<r�ڱ�-}�"�:	���)��)�b�����bG���|f�����`BR�(�}KA���{=�7tM*��EF%	��[&��bs�����)��ӅXC��+����ҪL6��W@ֱ)�zS"u@��.%�2�#�7u�ƚ�������S���Ʋ�Q Z�C��̙'��P���j6e�:�-�6�}�G��t�����V��Ϯ�;zv�c�O`��+�|VX�l�>Wpx�@�=�gF�1��Y*ƃ A��s�2��<�>dl���/��#�7����߆�[�놳�k`�c�}c)#��hT�T�2h#^�C�gly�j���H6��h�9ؓ)Pz��H�����Oy%��!{9��%���|�c#��18a��1�d#��BΕ�	߷d����`��'�$�|.~���rd�E�I���Z����	�Eȿ��2�P����9��Q�fݭ��Q%ȄE���`���S�دB�:À�D8��N�j2��i�__�y�AII�@oa�Ft��>�)2����H�n�?3�b�׭7Yo�0��H��x�=4s��i$���u]G����ցҏ���Gpz-���qMYi ��r""U�:ЌӨ)J�m���	2��"F�J��:�t�,8L�T�0���}N�\8�C ��1��j*�2����A����Kg�Z
X3:h�dmS`��luQ]��ӦE�����h@~.��#��L\���c(�(�a
4[a��\����G�[����
e���T��h�� N0m��4H�8�lp�N���	��(��y��6�ͨ�~�E�	̜v�)������66��B\�,t�	!��b#i��k	+Ѷ4|i���@o�wx<��xۨ5&,�#ۚ���rq�4��؍f14�H<�Ni����bD�ς:^]�]�b�:g���v�Q���C:��k��d���v�;�`��]=_}n������S�{��������	x�50yd��' |��uLI-������齜����9�ϳ�h�v�)aF���d�z�*����RgA����&93���"�V��5�m1� #+f@T��C��>�R�J�ƕ=��4��jp0��EP��3��(���x>`����P��'_���x�������+����>}��;�=��3�@�vw{�\㩍X`�4�G֚jԑ�2�c^0����P< ��Ԋ�9>@��@�>M1O�N3���e�K߉_á���(7Jz \d-�h2��m����c�4�oK���&�c�I��EM��QJW#
���s��6k�1
�����,�|�T�u-����=j���}���WV��xI��</��G&�1�S�}Ǳ�}k���5ՌU�YS�!���PC�	�\V���u�F*]r�tɨK��5N���PW�/6�,��_֤4�:�����)ʧ���``2d@ꠙ�:�z��d�O6j�Ĺ�L�g= %Q�kdTrs�ɤ`���y����r��������H!��Q����܇%�$�D ~0��I��O�Y�:��s�����lyDd�k>�?yCwB'e	��@���`�H�T��D�C |ȹsz�QK׭���(��:cF�N�E�6D"�	��}Y��S�5C􁾯1���_���׌0˚�%�� 3�^j�3�_\�J��"� u4��49�l�q��� ��l �=͠�l�C<���!�S(`�y?���)��ɢ��ި�鳂���]u��.[�r�-i4�$^Z�Ϻ�h�g+�L����P��{���k�lT/Y�2|Ǻ�[�c�]�JTk�玹�>��;���L�K�����)��\�L���ݎ%�\�j��?�甌WLT%SGmk��̕�K�&ImX&H�4�~g{�@K ��*�4�` ���ѣG噗^�	��:�/�q��{��9.H�ۢ�@��̬0F1�
��2�KO>��W;{Z�+����w���t�@PR�� 0��8C���{�_N�8!}}�Iu(c��5n�]���T�į5����0��Pd�b@*�����8�1��X
")�A�未AI 
��m�X����@�l@�[h���9`؟<���>T�(|�A��Lh6�A�#k�aN����)c�z��&Ř׀Ѡ^_i�A绽��1� +�Y}��'����]s���c���qo];�g1���u
�<�b�#����#"���拐55r�h4���K�馹=��jƵ��M�;��5�wj'���ΐ�9�^�\�{�R���2�,��Zf��N#a@��>M�u�!A'A3��BO�����
��F��F
&��t �f,S)I�W3#'\ ٨'��, O���rv7��+	SC�6�	`�c�� �<��C\ãIG3ąV]6�l�dר2�^k���^< ݵ�x�����N=��@+uϪ#����~&] da@k���H3�u͆���OW�S�W��D���6�����:u�}8}>bO�j��}����(5c�v)j�/ȱ�%YNN��_����k�30E�r��!���|/t����:@�R����|���" D,xv�#H�B�;!�<�R���P����F�pp$��X.)����^�a��}�z�#W�9�c���/ `(�U�:� ���٘x��:�FQ�1D.[���ԗ8F8� "0�M�J6
]��w
B�%�X�}����R'�"6��씕=Np ۵=�"�E�)
�r�U�6��3T�8��i�c���M���/~���&�3z���8��H��vQ�B9��e��i�=ٿ��n� �����G�Zm�ƈ⺑u���5~p {�T1����CCT��
�T���}�NM������F���ES4[����,s�Y�}���~�5����^\ާ�̓�O?!Ϲ�2���(���S,�W���P�	M�HG�-kv�#muf��TF{j����Pg���>�y��7�����lsw���������YZ� ��s���dol�(��dGb52㡍
�EYw����&٩�͓��H�fG����$c�aqYAO6�7(���Xy��'Ч��(����e��1)�&zj4K�҇�P�<���<,�Mi�}l,�#NY���cW�׻k��Kj<V��:H�%�KewX�{uL�́t"=��,�ؓ�:bu�Y,�i�4�W���;��E���6�5)d����m	1���J����b�+k����q$+=W����Y�<T'���fn ���͠F�ʇ�N�����֞8�O�:̾���|'�7���Q�n8���:k�?b9tiS"�O��3?� ��� KGNI�k���t�)��c�m��kD��5��Iٞ�j2� C?^֏h֭]_L���5	��Nv F4����4�����5�zU�<��6۲oeQ�uO7OjP��ϕ��4z���]^6���C�Y���}NL�:H8܊�`Ȕ����Xں�.;u��pi���.�� ��G�`�`��T��&Bߘ� !�3��f�A��}��MĲC�M��p�j�+Q�ؘ�GE���vJ�c]�H_�T }���o�CFK �C���( 7 �4�1S��I?j<6Շ��z�JP���R�Y;��U��o�yDp�8���ԁ
A� 0m��+Km�����N?~��"�KK��c���
���&Y�
HE�լ�$���'O��璘������o� Z��_YJEI����k�5#qow���KHzA)����Ϫ��.?ړ�X�k{o$���t�k�u��q E3��;$`mitd��)��e����t�o3i�|�:��ȼ�������p��c�{�z_��E����Lv{�yg4k]s ��$�����`�:CI6���:��A���������@_�+����-�>3f���M-R�J8()��Ǩ?�(�!���k�{pG��-+��A���=qRV�W$Q�9I=5`$��X���s���	�u�~]�"����Xև �f���-=��4��v����^ڑ@�s���B5�˭�&���N��! C����Mu:�f8�/Ͳ�z�w���@�#��T�k����� �K�&�bqH��pϓ�m޳86ed,%�3`�U����C�dK����O67��+����Ξe�엵�Uu�g��OD�֥��j'���ۥ�ò~蘍����'4�Ԡ3 Z
��	��$�~umE�V��g�'����w���d443�PN�Jۃ���:̺�����.
�x�v������5*հEB<AN6�NS3�t��$	��!˥~B<7<�UC��d�\���g@��h�-Jahg��&̽	d�/(��I�f��!i9����2Z�4g�Xǘ{��8��=�w6ͩ�,ld���91 c����w.`�֔qr#��&[S<݌�L�- 
�xn-{�H�J/��d}}{�`�d#�q)خ����8~P"�I$����� �Y�9�\�}�	d�dj���f�́��� �T���#ه�Ȗ��>�����<����l)��ӣ$�]7ղ:K��W]�9QC��.^',嚴��ޞ� }�ءF��z����J�xX}�p�\�_ȶ:�/�=+�.�ɂ(P�AAg�X��·��C����F̯No,�[N9{��Hz&�e���s������õ��!#T 4��i�9��#�b�@���f��[�� G����&mK�I(�Ey	�O@1b<ڠ���qX�#(Y������OȾ���N�  ��,��N�dA�� T������%��#`ゐ����g���M=o(S�!� c��J�=����(ooq�T�kI_��F��A��2�8�:�=$LFj|�CP�W�o%f�tcF.Z��-�ӏ4��A`���h ���YS�U�C���٥��j�w"0���.���k4E�e���	@�v�I����$!0�Q��-C9r���������`�_��!Q��SP���2=���x���֒:����Y���p����y��H��~�H+�d��!���o�뀈�t����Gi@��h���i��+��<�N>�1�ڤ~�$��L-�,�?R��q�"$��K�f�}�x |S3�CΒ�����x\�,Y�e�IbF��<���
AA���G��>�]9>56�1�9 p�G&Y�Q*D��G�g��T*n�t`�;w�P����/!���S�RǷ���a�Y��L|����5�N�9l���z�s�q�a���}-J�n�I_�|�,��8ν'n�/�}�5��_ [1����CqNP��*	K/0mi���:�5B���o��{����?���r\��w{g3�[MYZ^fo�СC����%�ڛ	K(��:�^����}+$K'�~eYbo��]&�6��Ƕ�ɒfCP�����8~�s�@r�_�;xX��9���P�@�i����{\����'0j��L`��#
t��4k�l��D�G@O/H�I!Ф�Ʀ�
�l�?�.zU͆���n����T^��z����@��#vow��U]#� �F�d��S�ME���l�i
 g�������Y����fe��"�\����Ki���e�/z��;�� ��AĐYV��f�k�Ɏ��{C��|�{Ӿ������$>�SJv��=O��D8�xY�ỳo�����F�d�)�m+n���ًj臂���쭁�M�,�'A���RPU�=@�����Cp!����p�c:���`6�Mܧ��%H��`�&)�l! ���?�k��=n�Չ��;��}�O���,�	E"��=�Af*C���0��bJ�=���u��!C5�JM�S�hԁP��"F�|S�!��F�8f���5F��$j���O��u� ?�H��.�� �C�,@x��/y�Ŝ��8ʻ��`���&�CX���IG����G�
Sf�S�O�	��s�kE���s��_5&��G��)�R��8{f��;7�R};עpζ�����ke��2�ަ<�9�6
�s
�-sB��>��S��pD�*Y$�AE�G-$Y�q{G�.���\�&�s7��1�����0���{�����Q�����&��cӠ��i5�ٶ���G��A��NhZ(�iF�h����f�L��=��^.G���'�ﻗ>G.?��ݺ�#�Ӎ�|��t�n?��i�����J�?	M�ԟ�)!Ć�,
�hN���}�2gk39qtU��
5"#̌����dHZ=�U� >V5��f��蹂6�h-�ȍ��xB`j��S��ܲY��ðt]ƛgfmB��EƂ�<��Q"��[]]�5��$}$ud3��0Ggi���ehP�&#�S�led`"[z�`;�L՘����Qg��:�RCN��ZdZ�Bi=%g�i&�IC]#�54&�0%�� hdpAC^/H�=G`��3J>N��-�K@����e)Ef��O|f��X���������0����J�C+���k���&��f��	i
Q�~e6FT�0�!�hj�`�C�I��陸=Us� ��FV��qQI�{ ���9��rt�tj��X�w��F�N�7~k*Z	Qߘ�.�?@!9u��PŪ��p�\���x���p�I�a9��z�(:�b�ecĝ5�[��G#j!Eh��6A~�2t�۔���ɲ��U�nu�^Y�u���5չYY���*(��#w���ԥʷ/�uA�U�U:^�����J� �a��}���d9��V��95��	&:�W`.0ҡ�]�,�
gLR �r���Q����M��dD��]^^%Q�/�⇞��g~J.��w����8�b���ٛ��#D���:��.˨�>��:1�0���G�f�l�ܖ,�5��M�n�ȵ/�O-W8f}�vD�����8$�QK�`�X��$R�5k���Z�ĕ0*E�*%�B
�N߈"�p�fQ�@�ZRH��R JD�ct(�$�VR���2u`�'S3<0�d7r*:����C��l�HR�`���9�99�M�畦��p��J�!zng�P�8>�
�b�@\F��?p,A����=s�� "�f �e��3�bL#M`�eN�I�;�c����=Δ�t	 ��g�;@�RP�`�$48�-��@��r�)�\T��L3�+&z�> �}�V�##��e;2��#�(��e6��Qt�@��rJ�����6�����5��`�S[�B��F�ꄢ�G�j��	9� ����M������2���K��sn ^`�&�K�n����t�}���e����pA
��_��Q�)K�Q��sU���:�Ӟ9*:Rz�� ���)m��!+[���޾��w�ϥ� ��Mޢ*���&�~�C����ܕ�q� ľ�]y���YH��L��`��T8zF,�Sв2���9���r4�����+�� �=ڿ����g�,A��s��>����g��;�9��#�Ϡ�DEq8}��+��������}gk�ߟ;�(�;;t���QN����h L/��A���⥗]E�d��d����:��\�� ������`C��@�q�U��W�	��)4Pp@��Y^��U�0'�cC߻I��O�n`��@C��&KK�p$�a/�!��8k��#�0at�z�q���fU�%�؄�ۚ��(��Q�B��â�F�A&'=g������$�L���f����'��;<�Vr&AJPcy��u��A��\!�g�)`y.��ɹn�MN��AR�2�1����P�)F�S
���=	H��<����K�KŐ�	D���ӡ��=�"�˙)�0B����9{_ߕ$���W΂eV���P�,dB���l�ٔ|�1����Q�>R�^��,;�H�u�Q�Y����7F�l�@���E��~����"X�87e�DJTJ\(6�u�BND5dߠ��4��3�5zb�<�[c�C�A�qJ���م.�-��� =hn�[XY��VIڏ�aϗ���,�)$��Yf������F����i�P&�'n����;Ϯ��;�[f�6>f�cU:�dh�}L�&���H��\������9�۞!��D=�W9^�9���e���Ži�]�[��]aׇ��l$ {��e��"%�F�"Gs
[��yd3�$��g;���~tG����:�\��r��m���8����{����]�Av��z65,+�i��p_z����@VV��D�٣��l �R�5��C��DcJRې��7�L]aYX�Q'��Y:��lNA霽a���
�:
˽�1��@ƚ�N�03�Bb����)K�(��R�! U#f��G�iz!�/%��+#;t&e49=����A��*�z������3��>�(�"�u�EM�f��,�K!o��l��̶<�1[�0�-k�yf=Q��dd��g��( �v)!,���B��h's�`x���E�m푑��!N�9Όl2�N5��Հ*���#����)��:c�1��\{?T����o#'4��7iի$�>���I��K���LU&�����U�D�^6Ȃ~@����~��3��%*A�G�1�0�T�;��9pn�A�(���$�a���z��?��Aa�fj����̬p��I���[ꔷ�ܕi��sf��*A��F��>���4���}O��z��"��uB�����>��̦,	�dKdY^e�8̉;@Ra�q8d^�����q��nT�2M��R;7�]�`�Ì�8GC0�e�ei;gߞ��r��Ʌ�� سЂ��3��_�ئ�fUJ
�ͪ	�_V>�� K�Vg��2�mku��?��cC�h��62���j��0�I�یeue���E7��7�<.x�{�Wn��'n���~���{�u�K��'���'[�6���p���No�k���0��S>���,�v�5ٙB�c ��\I���CL��W�_����2F9H7h=�g4 �H�0����i%��~j��$��-!{0#�&r^�L�=ѿo$ �����YV��|8��؅�4@IXl��6u�\�,f� w�YFN�r��g����.cyJ5���A�>�����,5�x݅�� [hj(�[�F�w�Պ�1KCz�5A0���]Ru�9�b��FS���~괚��Ҍ2���k��Hd7:��[�t"pz���YZ���n���E0�%�D�}˄���R�9e�9�l F�:-�Dd���ν2�g�Y�g��h�Cd�
��a���a`2�\1�� Q�>�]`�DT[<qlZ�+`��$-��X��������y�Ey�8�� ���I	`B{��܄N�[u!t٭e���9�b��� i��.�2q>X���&{ݱS���'>��N��!t��W�g��N�{՞2��S� �F�W�d��dvne9���� ��+�&o��RQ�:��y����{�Θ��V=q���ר�g�ꐵDy|iyQ���{�N9����@`B[�0�74 %���ӱ�o���r[�A�?|���x���x\��G7n�����w�q�j'�?��]hO:c`T�>U�P6��f't���ٶ���Ơ�ӌ+���<&z�F�o���z�a���C6�_�<�������s��*0���K��!9�$A��,WX�<�=�^�8�ss���9ba C��!/�ÍM\~^���M����(�|���y�HjD�z�W��`�2S����ʿzst#c��)u�)ڐ�{煍�v�dT朜����y�^�}^.��z"匦�;�&9�
�l��:;�'g2��?��Q�q�J��s�feJ���,�z.cs�!I)��j�&���pC�������5�]���y�~��3gI���e5q�E+=ۓc���P��3����&���;Ή��gY��
����wc3�K���y1��8K��8}��@`�?�|�B���1��ݞ�V({��ܳS����ܲ�k ��	�N�˃rd��Vnlwn��4�q�s��wy�Rrn?ՆLK����G@\�o�!����'ZQz^O<�V^�F���>� *����j�K���=�si�d%�1�Ϊ��x��wr���]w�=��������/yF@卭�LF�� [	|��3kqN'��(�R�5��:F_��N��1�l�Pڝ����bN35�{x�rZi�f��C��N?gY���=�rp^aF�(�}ߡ(�2{e�S��?o���(����P�$�:�u�3����7I�)�A�^� y�����(��Qڤn1�?��ê��n1e)j��B��
���UC�f����z���^�s�����ū�yY����)9�_�d}�Q�Ѽ��QXhhe�y)�*<;_�A�J�v[�3�^C�{ޔ�t���Zx��2�
�V����*�9����x֗+�}'+������=�$Q��ln�f���@r�^"��>/�W8� A�Xf[E�#�a�l|Ԣ�;p��LJ8�7�I���=K��Q>#R����gFs*����>�g8�bZЙ؞Ꮆ`	���J�Y��C"��z�\_@��	����v��=a��A�;2�Tmqk���l
؂�<�Zv;���I����֤ړ��$�8wmu��=�s擔T�Q=����c<�*�q~�Ɏb�@��b�X:��67���$��}��x�s����/ߔ���x�qճ���O~�3������.���(�%.�d))��`Z�>���3���`�0��Ӡvm����Aco���E���<
��o�Y���dş��i�(߲�³e�ˉ|����?��ܺe���g,SY6��~i�oD�ee�ҹ;�n8��y>��Ν����V��*P�q?����]6_����J��e��d���-#��.�����3=�3�r^9�H��C@y�Md��]���݊R��VH�ϱ(\Vl�O_��K=������ys������0.��<��R�#w��sg�*G��~�����W� +1�6W���lp��%��Yu�+Q�U0Ŋ�Wq!��ܛ�(���ݾ%QH��Q�rfχ������Z:�¯�"K�9����Rl���L^12O��1F1�;���6� ��' ̲r�`�r��K��������Xp4�C
�H����Oa3�l��-~�נ�3���E�@㔻�unh���ƬO\T��=e��|�l�3i5���
S�2V�R���<�"$y��]��5�aN�e�@N]u�X\����ߑ����+�>.:^w�|�M���[���νh���E���`��ȴ0���{��X�"l��j>$����Q�����0\C��	F�@�W���tse�y^�.��.�/���~m|Ґ�~QV>���b�.��B����Q���L�v�<���7��2K��eZP��{�[�Ye	�e���u3�0�R�oh�}�벉�(3z�@maL���J1F�.S�Ls�M��eaT��\��'��ݓb&)��Qq�!s{��Xf#E�S,G;P�(ת(��b���(���.3���.�������9}�9 �Ci	�C���dS���4��s��C�.�*H�$v�y��^��q���!tc�*�H� ߭'Wn�i:!P��w���*H��������:�ѡ�w{��=�BJ���2�s�%q�?W�(��
OTTȴ� ����t�V,�Ǚv�9f�����+�s}|� 9�\��v��E;��6Aͦ�Jb�(p�W�D�����@��n�(G�b�� cy��6G{�R�@/��7�T�K��d&��O�s��]����رc<'$���I�B����&7�bJ��l�����lwaU.���;�~�e������={�88�1���g��rQ��-� yGD�ɦ��~�1P�YH�zA�|��H�F����q��ƕ�/��_����AF�����G�*dΐ��Y��r�);*:)�
���
��򌡧$�%��3C��#�3��YDC�Y���Y��yU^��=M�s����Xeӣ�)����5;���ЀD��)�1�b\�E�E�Ww����ʉWT}�y'�Y�㜭�����J�e����2G4R8Jǒh�~o&���>�2����q����%�O�YVGU��� �EQ�Uy�m���z�  ��IDAT%����\v<�������\y>�k��i���TS e ��U8.����6�l��\�\�]nFRq΁-��=�UʶK����E��#$Ș���C2���5��<�����BA�V�73�q_##��I���ρ���a�M�=���t�5:*��V~ #@ܿY-Gr��D�Z�R�[d�t���`�Y"ά�Pr?��ZR�y�Z�T�5�w{�J�ϱS�5&HRR� $�K)�v:�����U����D%�tL��)�0&�טj�+pÃ�jkgO�����{A����z\s�5����?��w�}�{���JY\X���m��3U�a�9�^I�������	�OY}Uh� �Z�Fq8�<N�����ѧ���e �ӿ�5����KY�+��=���k1�S���Y�_eeR8T��g�*��F&f'k�?�H�^�&�I�h����s.���yV}��ܒh�L̝1��������~5G+�c3<\�xJ�E�׳,AE4�E�3 at��n= pE��O�,3�r�ś�x�x�b�_l�H �#˾�#+3��s��`��o���g��h�ع���fߡ�m�C� ͷ3أ� e�Ue���qw�;什�e���;�9�zB��2c�J��z�9�����$u���(p��Q-��m�����[b�m�c�5�Uov��9��Q�mk�X�,;D+�]�Z��fы��Oe�y:6�'���e�y���m:~ �9�>N��;5Ǉ��_�x��_2�#�M��3-�*~J�j�\`(MIj�sլ6����s�܀� �����ƙ���ӍX�'�� �yn f�kj� .��ݒ���XB
1��O_R�@����)��n��Wo�/��z�����;e��Y�7M�de��$��x�#՞n�вD+U�2� b��z�a=�1F��f�l�}����ʃ�8�<���rFO�tx~dD��U"'KTf��S���1��>Ӎ��?�O��!ՠ H��q�a�o��gN��W��SϽ:'�	fY��[�0��Jn♱*_���H�w.����zA1�,�#����u�HP�=A������љ��=;�zD[�	�`3�yyoq?]�3�N-צZ++#��R�l��� �}P?�fS�=���ue��xv����F`��;/�.ISp�3?���oE~E&aI��>#�}�͛�y��Nٞ���<��+,k.{Ķ7l=����2��v��Oթ%��%��m���l��}�e��w�~h�擌��/,`�dS{	���@�z�l��l~�7��GcUY���'��^����Ԁ,5j�b�&s՝��.F�Цj�=E������v�YE��$�k%n t\���:�K�;�R�����@���.�Q����9���v���)���hw A�'p�c�����48g�5xP��������PZk�;�s�����x��8r��O>���9r,�5�9����(#I���0�����F��dL��zC�T4��D:(��ΖF�]���v��PM��ey��eY����2������ɖ��Oy_�*_fU�T���|�D3�y��TiQ���>�ޔF��/�19%����5��XY��A��9?9��6>��w L�\gwfF�Y�T?/A3�
�c�֙��G�Ȋ�;/�K��Rz=M&�ˁ6���ȌƩ�D�-vF�4�p�|O�D����u+s*C����Og��� ˵�w�֋ˍ"��zѸ'�������A0�h�_U�����D�j ��9.|RTR�N����~?M�9�[�V]U��h#������AT��Dv �T�r<ʐ��zu����7�α�=̵$�0�y|�2�9�rO�X��}˺I��(2�J�M����#?��-zu�h�[�9-���M{���l��g=V�Y�۾��8��M���d�f�I�"�=$�?���}�I���$Y)
����6��k,��G��_{�1i�����yM�,H��	2T��"d�7���{�ը��P�Ig!����\�U0��b�%���,v�i���u�uO���k���� �b�
9�6b����/6��EA �\Tv���/}�K?�G��uc�nyqI�=5;}jJƎ�f�'���s`o U�	Ӣ��Y!TrB�e ��h�\�p���;+���\�+�RLf��U�Ӂ(lp�H�Y@sY��@&~�QzFLPf}Π��'Sf>�m@����9M��8˗�f��i >�3�iح�[��0���R5C�zx���߳�X6�gVR�o��kl�i�mN���h���N8:�C5b����`"��6��4��j��%|n���,����'Kښ�E��~�߁Q\�u8s(�����?��N��Yf���%&;��0�4�.�(�����
� ���:�qY�50R����a��$g`�J2Ω{��W�de�yn�<�ys�Aa#i�ʬNd<����F�'��-@� �D�X���=���!+޿7��
Ǎ�엳�Cq�_E�X?�ٳ�.�*�Q\KɤV6��V�Q#u�p�u���E�����L��ԕ�JW����������{�%�(�qǝ_�e��Y�:¬+�g���J��&P!n����'�˟)_u�5���epv�>�7�(���hA�u�����믗��KS��h�IX���]@W�6��h��]|��v g���n�v�m�,�E��Lt��ҟ�U���k
:rh��Z����;6���$Ĉ;3׎�I�~������K�����fu��3�;���ۣD`�$�"��Uɧ0BS)qą3^idz�h}L�#2�	��%뀵���L]��j�5[�g%����<�<��́��(�c��\�{����sr}.h��)�o�H�N�e�j�B�J��XMX O5��d�>.����7�Q6�,~��,�pb��D��}Ą�S��I�4��qc *�a����X���A8��9#Y����ׂB���\C���Z��J����8
Eq�	�7q�!��/��Ը��^đ�x�Q�e���|�U����|��<D���X�0����P���� �I0�0~a�8�f����MC/����'#�`�N#��N�{�U�kϜ֔`���L������`�ZCsY2���%��<�k!�������VL�Z��t�0hÚ�I��L˽V)�h��D���@/��+��k�*F�}����2:ދ��3@S(371dү���|���ܞ}ɥrdmM��|̮x��PUhՕZ�X�\�|��$nY`�#'��^���_��?q��t�Y2�i@�e����x.�����o}�-�t�O}�3�o}?�WU��Q?V3����o�?q�W�����Q��
Vؤ�֫lw �9JQ��n��L�1�0J�6|��gԣ��7%,�8
���;.:���e7<|�������o��-k�7Ј3��ş�7څ��%���D�Sd���M�G�F�Yo��f�0�3t��"�+ź�Y��A	]߈����]��b��r'C7+\#��]&N�`:W�s4�iR��ٛt�S���6'��,�s��$x�k�L�~��S�+�\S3��s�?�����ڟ������W�4f���⠡�rZf8�w�ѐc��h�E	׌l��djN17��i�-/b��	L��ۋKv���������VD-.2���1f��{\M��J�Q��j:���I����!e�9�Ǉ�+l�Ӿg���k���s�����y�Ĉ �tZ����qISz}�-��D&�\F7�?���Y����뵦�D`�2?@a@
�eT�\��}��m�t��!�-xE�����3'������No�LP�l�=� D2��J���p2��Kb ˋr�+n��z�|�����l:8+0�P��Ŝ$���>S��f�Ìt��nG�֗�[n��=,���㲲�h��}�@��V�%q�e�&]�o��o�3g��m�ݦ���[[�c#j���ԗ��6֨��[닗N��2Ynԝ0Dx&S�}��g���N��rTYqܦ�f���=p���!�b�mҢ���v��{�x�㦯�����G>��e	nұl<rZ����R���N�K���|�9���ʔ`tB����d����.�̍��D*&i� r���������F��U���ƾ?3J�r�@����?ʦf�WI[XT��FȬ�����,��`�0�"�]��)�Y��
O3�q�8���5�I��X8�3��~��*2��T����Q���(��|vß�}�B�l��2��i�:���WQ�(_Gɻ܂��Dc`� t����`
&\Ʃ��${��R�83�&���g������r�����ʵ��j>%aU��;�(�"L�}�u&Ƥ��J����,j��sF�@�K܊%�8�V&'U�ó�
�05�eՇ�`��_D�f�ӌ�qj��q�b�`��"�G���	�9c��G��:��| :[�2�3���vK$�=U��J	
��$�L_(���D�o�n#��w�e�~�����𫮗�֞��ϾC�zu}@gӁ�)�Ñ, h+��5!p*�p{�+K˫�7�I>����f͇� LQ�:m�9SVg�$֠ϋk�}�<�Ѓ��������ԣ��2/��k��Y1r�.�UMP��KPu���)�x��ލ�;��Yn-ҮS|f���h�:5�S��(�t��<��}:3�{��l���r��?sؿ�����3{;r��?'�ӏ� (2�\+�3w=O�=�W!�����@֕�� ��Q���#� �6Kg��9��qE�+��.�����2Zz>��(OsN �|)��~!y�r1(}GFB/�\�L�	8JPS�L4-4#�v�._�u���W<[R����L6q_V���s����ߗ?�5�\Q�v���!W9&�������rҲ��8:Ð9C@ c��'I�����E�ǼF�$�nеN��i��(��vu��8�CZ���ey#���&FD�bO��$���C��.��1��*�	N`u���sߣ�4* �~��Y���E��ɕ��.Q\�4@�z�R�)K�X���O�8��!�g��ʚL�u� �y���Q�� .dP�$n�equU.������s�ao����?����3�`��c��c�h�^0�C��].t��
��K��Zߜ2z��`$���ߔ�C? �^�L"�����mrX�)Fbp�z;�u8�t�����\e	a *I��7��o�G}D~�w~��=�Tת�9��B9|�t5����w|������|�C��* н���R � �(�`M2��31cK�#�`P�-f���g��D �L�a`����1�1c���> /��\^�>1ޏ� ���lEP�j�E0O�QJB�u�]t���н��5��]�%�j�4���  F��n|�d��{eI�"�jF��J��u'��"�(�g��p<�d��Y� ��'f��4��]Ȥl�ȑ!�#
ۗ��%.+��^B����0 P�m%X}Ȣ�e\��Y�m�Y�Q��S���a��ѱ���6K�r��)� 
�VgFS4��F=�8������fX]��w�iitg������Z5:¿	�,��T�"W2ͨ�k�624uq�NMG5�����@���Z�E�i-,:zg�,p�@m�a/��B	�"���"���"��l�ê��B�Yϭtᬊ1�1e��U�#�Hu�X�M�zΏ~5��ң� T3˙�+��O�����=zT�5[?�G�����(�U�+˴e��u:�8�?�}j:��k����j�޿O��_�{�Ov�{���&����5�Y�y�&�h�?��X)ޞ)�w�6W��#�\��VE����= tA` #(XV`�d�B�7%PG�����>�`O�����)v��Z�a���IR����s4�C\���,��ɫ����Ï�o��~����4�h�9e�=�j�����th�;{��W�d������Wj���aGV�]I�c{P<�4���[��?#�����ˍ�*QJ� �F��%f!'ZzW�b<|<!e%�.���"uyZ�=;ɓ���9I}�M��Aҋ=ދ�?}���'���@ �հ��83A�L���H0L�=g摖y�d�.*� W``�~�A�#���E�#&F�F�7�yD�p�a9�.�4}iv:�lkydeLW.�빡t��5���ˠ�ӇS,��K��d~6!��K�,R��eޕ�M���X�EC�iZ�,U!���:�z}E3�-'}]��$aNc��5i6jd�����O��S� �F��Q�J�Š~��׎kB�%n8O����8`��@_��\��w�#�}�9vTt���+&��4���us�(�����}L�{�f;���x�h6Җ���o�����b,=��� ��mUʇ?!"y*O�~L��	-�QE�u��2���F0�k����3���P+�'�����HӠ��!d�G]p�T+�N�)KKVR���c�BI6��H�&q���Z�4��2p��'Ƙ�vR���������}���|��F��4������|�O>*�z���,�o������Iu��Rf\�Orc~�#_c?���*c�8��!S�L� =�D�A�/��s�j�]����2V���|qiɀg���XY����ż�Q�nBɚ��bs�2�(��ri�by��ߨ��P~�n� G��BC��P�)�#]������x��tu�W��."��x��#�@� �cyy��O+�[�pd-�M��lt��mf;$EiJ�k<Ϭ<y6�nHp�=x8c8f�H|�I�4>g�^l�GA%II8��;���f�U����z�n�-�n�iNO��9.:�� ^I-p�~�ץ1ܕ��Ӏ�&�L��F	ܫ�˽�	Q!z��5���=�`K7��+�9J�0�qy���h	"f,4k��z�k���LL���޶���1(�\d�俒��� ���Z|Yҿ����it�踣Y6���P'j���u#d
�t��^� �F�[jH�Db�n�p���/IT�Js�&C}��\�b�)�ͳ�?�S9��f<���F�7������_����A6�N���k��_|ܘ�|s̸&d����Dn|�Ke��1:�t��n�59�F�_����+�:y _������ч4Siʁد��3���~ӷ|�<������R���k��n1#�
�J�������H�Nl;fQp�<���u5�q���}��S#�{�];n����#XM�d�g���_�My�O�� ;��r��F_#Hu:τ�u�����	�?��+Ca3M�k�3�h���~?4f1�	�ܣT���m�.-�4��������ў�k�0�>����z/"�Ud�8,p�\z���Ⱦ���/
��6�C��u�'��a͎��%��9u���L��k`�'��uQS��[���mr�]� ׿�i��Q�D�>r�Ü[mu����a9u�eƲ��i8�P{,w~���?��cuuf/x����� �#kz)cY��Ӻ�V5���?�C��:��m?&�nK���r���t�\���?�����Ç�4�y�=���Q1@{����G��^H��z�5�w1��.����f��ّ�x��j�Aq��pK�Y�6G|Vڍ�����@�U��M����]��ృ$��2��9`|�]�W�ʡ�"u4�4��9�S��o��A�kd�"�q�s+���24�7 b�jK�x��ZV� �fa�_�{���� �L��	p@O��ɢ-+��k�gj&7wwj@9�'�q���3G�G�͈j榡$�3u�z����9��IF������Q�	�ptS6bA��� ���=u  u`�Qr�<����WĆo������F<8o�r���^Ї���
�z��k�nU8i�����Tg���.�nW��9��IZ��_�J�R��J�f�� %*d�����:�z�ô/�!BK߿�q�@?�5�Y�4c<yN~�?��V�W~���Y^`������������W}��8x�k���:g���~H�V��p8��3���m���w���o�Q�k	g{Q�\�5$j��<�/�G�����W�o_�F����f�[��_���K�$ߕ}��@?�I�l��l�:#��^�>u.�|�7������^�^`*3��t�����-��	25��	ztM�RǶ��jY�&� eY��P����M��OlL��U����iֽ�f��}Dvu/TG�J�f��@��W���L{F����$���s�=u�<t�]XĲ��q�G��Y����?��e��K�����ˡK�Q���������9�]!?��w����'k���|�����"�V��,�>��
�{rngC��-˫t�k.�D�d�Ց,���ǎ��C��8Gr龓�J��o�_��S�Nɮf�>��<�W˿����{z]������w�������d��4t�~���ʒ
_u�_�ߌ䁿�C���_�gŗ�~���ҡ���mK_��_��wɛ��Mr����ht$��ߑ_z�<v�I9���}n��I�'�;ĵ�	���l������x=��z�k�ޣ�k��k;�2ل���xW�^����_�������W��:A8t"t�b��>))]�\��Y�x���`����p��x���x�f�QI�������A��dQ�0hʌy�Ҕ�G�%����y��娒~�JԒ�s{j�����|�t��'X������tG�~�o[Xd���<�)�P���>����+�Ob'����{d����R�1�A���{R��L��c5
`�aI2�����c��t<d_��Qu��-(3�C��X	J�j�0�[#��v�X�#�������ͶZ��x�["萔e�T/mO3�Y�zW��C^���1�D�z(+����;r���_�u��YWț5h�-���i�{��׷J>�����~��/7.g]���<�YWj�5�I�ٸ����s���>��w�S��3r˷�K}Jƃ� lj"��O��_�
��[^�k=�v7IҀ2�+_w�f�S��?�Ky�Kn�����ވ@���mK��6=��%M5�}?��SZ�;M%N9S�@�&����-���;��^��TS������Iٿ��k���OJ�=��ş�79�q�\y�$e2R���[W6�<C	Jd�yݷ���d�Ҷ6�۷ʿ���h�p߃ȓg�������7�A=B*�о�?���/.�ZwE677�/�ǟț�����3�K]��ÿ��r��/�g��B�z������}���%7�(W]u��s���_~��F����5����ş�y�s�+_�ʯ���wR����|�O���Pg|�yW���R�Z�h=�
��|�_��:�%�� �2@�u��W���z!���9����Ӻ~�-?*ϻ��A��{�w���������7�NoS>�G�/?���<�yϓ��M3�uz��?�g��:i,td�N��D��O��\v�Y}"��ٟ��5{ٍ/a�7�F���y���O�]���?�V�>�-u�#�c}DJs�,�Ƣ��zͦu�.��~�+���;��OJW�0�&��Pj��w�N1��$Ҡ���My��{y���C2RG�m]��)Q�2�m��E�
5\��BD�u!�$D9��*��8}͒f�p�,W��X{	�B�(h�����g>k��C��pL��<d��z�^β5�8;TI
�v#qP�=vo��#�@�����9�k(١�J"�xHͻ2����ӂ=%8I(ǀd��kB���-}�:����T�2Їfk2�^��X��)��جk>���D��7�y�2!{8��f5�-AÇ(wm�+#������o��D5�%�s�,��n�æ�m+��f�}ϑ~������X�V��4g=�1 fj�Qbm���K0S�g4`sf{���o>�I���������H��,,�7���r�=��C��G�])Ya_`����^�H���}�<�9W���-]���������L`����P���2��s�3�h�׵�����(?�o~@�����k_�"����qj!�É��.�I����2!*��#YY^��S3BdzK�T���+�ӏ����M|��>y���}P���?!�r��q9�����?_N��zIj��6v�����o�w?�u��m�w�؏�[~��r���5��������s�o�.u���}��?�S����M�ɟ~��ܽ�G~Xn��������o�d�|@��K�\����WM��$����$o~��军_�s~ε�� �2��=�k��\�M"Xc� ���7��+�` zr}]Nk���D~���d�Xz��}`?v":�{�G�j����Z��>�z�I'rN�Ƿ��;��ӧee���y�	y�{�+߫�~͋n���])t���8)����?�?*/��zYV��η��@�QoOF�;�>NV�K/����Dǡ�,��������뽹�� ?�#oU�'��X�@��k0�{q�חH�ݚ�ö:V����8�:���4P��5�LpCFXKu2_�қdU�O��t6�@�+���g�< � �4vk{C����d��qy����ۇ���T� �[�ƥJ�[P3�)�*����'��ي��C���}VA���{�' n贝� h�����Tl2�; 9Z9ϱ݅�L�cC�l�+G� �@��H�%jwX9���d�4����x��#�R_7���)��
 M�n���U��M_��h#�*R���/ 
�{YB��@.A֧�2U�� ��*����f��{�ᡲ���f���uBat����YQ�����~(�0���Ɛ���Ld�a����.-v%�M���9}`������}.�F��`�態�G����c�=�$;�k�}ﭜC�0=9�(��"
H�@$���d���y`xaLp �1IH	�B9����=3���rݺu��ϭ��ߓ߿����>��t��u��>�9{��ͤ_���R�pc�}x�>\�⋑�M�F`�2��GR���%(�}�_�ʥ""1P�,z�3ڷ��e�UZ�B5����vaA/}�ˑ��r] W&�D&�lt~��pe��F�QJ��{�VVg�	�|Q���V,Á�q�%iz�
궊�0�*�#Z��o7~����jQ�[_ s���k���a��tݛ���9睋��ڊw
HZ1r�N;��B�m:��z0���?�1.8k�}��5� �x�+_���)l���x�i'�b0ۋW\q%N�	{"7�x<�K^�Re�͚�IKF��_ߏm�6�_�ip����oVn`�Y�Z����(y�yϯ�p�E�aکX�|6�x�J=[�����zO�?i=��^�ö�N�E�m Y� �U�u�������w4S载Y���t\�W�����2����}{���V�#"�?3�#�1Y���'����Oـ�o�C�,�ͣ0�?~��8thq�N�PL�qx��sr�1 � l�0?]Bvx@��:�׿�J^�Ρh\�-C��"�\��a�1���P�m�vn�y M Rф�hK�i�lW��U��eD��in�zI�\nq�g�B_��2^�Wc`�|��C��)y}M/(�O���[��<Tcm	ԌY:��V>_�#-�홏,�:��2�gq[G#�*`A�C��{@�+E͸�Y��`�%��v��:�6����{�i�]�\� P���gճ�cD�I]�S�{^��q�J�헽�-�q��.��0lS�[M�^�=�T�T#����$;���F{LK�0�ik&���VBAn��dF��|F$��0�� u�QC�Q�Dߎ��Pp�[W5�Y����L/��b�l�V���=�\;�Ip�'�a����Ƣz,LC����s��`er[�8�cA�C}���^�S�F�]�k�`��w��|�a4]}m+����+�ۣ�x��)A�c�d�r|�w= l�tN���6\{���t�U�f���~70J�ÿ}Hӛ/��2e�f�7����h�vXXTO�ퟷ�^�M@���j
�>�%�X�j�:���LO	b�W,�*nϐO���(��)�HT΁�옪B�RZoH�۟�����|߼�+8�ҋ�I�-�
 �X�n���҂w��$�!��{��	`М�T����0�d�L�9��Yi�D���C����q/�a�/���^��~p+�����(pL@k��U��W <ԣ�U{>ի����;�rW'�~J'�Uଠ�T�ZD�֠f[K:aR�l"�X2�K/\��7jZ�U����/tl�R�V���Ԋ~yMv�[�l�?~�s���7`J��P۸,��cmhA���jr߳r]"[|��Go�ox��]�����������k���gl��s�<2�+�9���L��� v�م�[6c�V����)H �����]��G��zE���c�-ޓ1۫��N!>���EV���F��,.��
��af�EI����Vj��S��@ �4E3$pbA&(Z��&U�a;�i�Ҝ��0X|�����ܪ0�Vӫ�g���1�Dh��Ǧ�3֛���L�Q�/h�������9��C̟=;F�%��7=̖Z#��S�����my[�	1�������S8�������wv�É:���ñ�m؇W2O�I�e��I�w�=��.�zR�
:x"	\���[4�v��
��I�,�2N�G�Fk�{�l->��/Ӫ*�Ϣ���=�������u��#�u��Ý�GJ�̀�/�5���Q�ʷdⰽV2vyO�\Ԣ��LR���s�^q�����������>���}:0Hu�Y��B�I� �j�H(����_��	�e��	 �Z<���?�)�n
;�	k�����l�!�1u-��󲫮��SN���ʄZ��5m�X��`�%F��r)��2��Ja'a���)�  �g�֬;I&�(������,r�19΢\��/��Y��0���\X�ip�u-��kN:E��4<|��8����Z�Ut�B9�@T>�S�å�h �,�jW�r��5�_�ª/�r���q���{>�?������O']��O�H�oto{�;���Ž���͏��}���>��ϫ�o"����������RP�8� �gK�H�.�!7��ɵ�j֐�Ia.����n�����^�K�'�%���\sC��/,����y�h�ZQ*���}��G��G��O`��5���˳�W{���#j.B������{����L_z���j�X&�\� �s%|r�#����S�3��[-c�)��$���0�r�6��cLw���K\���:.���.�k��E�Y.��"�ȹ;��i����+R��IPdԩ.�;H��`{KH�L뷜�(����.#����sڙ�BIS��)�q��a �Xq,�[�Br^��������ͨ>�uܙ�].a��v
��Ь�f6���L�s�rlzE���v�|�U��O�Jvz�ev`�J���:�#!�z�d���2��۸�=�����o~
'������͎URR�}F����U{6`F��ӳ�z�����Lo��`ݖ<0��Y�e{Fi�ܤqNVH�����$�50��CզD�m�PS�)��k�k���sK{4s� ���a��%���Т"M3�@GP�K�o̎��lC&΅�%��ͣ��-���U����yp�@���i�Pc�u[���;L�OONa���([Nd�d����d2�!��̶'�Ľ�I b���ڕ+�f�j���ߏ�L�u�LȤ�vPeц	S�3�>	2"
b���"p6��	�����Nbh�_3`5 �4��<���x�$�d�:��;�M�JT�D峪r�(��I�Nv�3o��9Yc��{v���{w! ���?�[֯�,��z��t&�k�a)�0��/y�8���.�z�����<�	��"S����/�R"��P�����*(:4. 0�����/�b�m>��)�����my,���[p��oS��@ ��#a�N3rE��j{���J55�pU�!- qdf
��������M���= ����j����N&8_������/���sT�%�w�+��m�ܪ}�gl:]���CGp�=��uo�F���E"��ܣ���lظ^��;�|
_��?��5w�7(W���M�=�l�Fg��Uo|#��կ��'��5�}�
�}��0#�b= �"%���^o>A�~�=�������E�c�� >��1,C����T0ӊa��%�hV�h�j,ڴ_���bY�5�&L��;ecr�zĚf�4�az�\ˮjM�fG�@�y���޼�6���^�J0�gJ�ٖeq'�b�f��/�<iZ��A�Q�;*Ik�m�kO�R��܎[[�!P���ذ�r�^�g�ٔ{���P��낫^����oq"�.������`f�VhQK�JF��ou=��c$�['9Vw��ǫ�˦'�h	�Ζ
Z4��E����Y���~���i��Y���	���Ɨt��y���T���G5m�@�X%#�|o&��+u���D�x*ג��@�g=�̈����R��(-(,������L����,�h�Q�ϗ�4)��5E&�/~����I#�J̏�L$NޠVfq�9afM�I�Ӑϝ��1&Alh�Fe���4|>]�Ղ��O�UZ��Īk[	Ơ�EV��r׽w�
�\c2�%�&{T%),��w�LN�ɧn@-��9�����P˔��E:,2���t��W�N�����~WC�>I�\/�_�.|��x�K^�?����;?����W�&ݭ4K�{�A�3���݊իW��F0�BQ�����fq�{ޥ׍�r�J	k �V5z�2s!�(��m��=��
����
ZP1�T^֜@�?KX`��'eQ>�od�\�b|�_P=�E�������.����/Ӣ#��w*�D܋3���H��0X� "�M��tN�"	-	�jXu�r����O�����e˖iF ��-�~;B}��8��i�7��M��߾�k�%	j�ڲ]�2��&�-���x������'���}�߄_���Y��%	"N=�,5U��^ϭ#�K�w�?��V|�G?�@(��]�:�⚫5�P�fq�.�!�}�$@���ˀ����Y�^��a|�cF��"�"{W�R�i��ӵ"6^p6��ی�|��K�1 �HB��KC*2��L	h�Z�h;��+�9i��QeL�y&��v�7�*cf"���V)�DgF��_[�ѿ�K�,�Q�4�k�650L�ҙ��r�H��F�!��~p�iz����V��m��I� ���ܳ����W\�g6�|t���e���2�V[���MmYUv�B�s����&p�j�Ƕ���!��	���ziM��|�[�a�M��B�<��rE��znA{m����`�y��-7��ʕ���C�M��=rYa�	38>~Pې\�!�����L��[�db@&.aT��+�ˇ�)3
�T�e�t��f�g���8�71ӥ*k�3����_�/}�3X�d%.�+�p�w�BS��J����İP�[HS�U����1;7�83�P��m��j%����*Œ6��	���Q��߉���_Ogp�L�K�1;3#�_�-[�o݊7^̘�E�*� ��l_�}����Vd����3X-�P�i`�PV����n��.`�I�Q��f�0�H<����JL���w���ߢ�(�8}�22������P��_�~���aÆ�V�u띘/�q���b�ikP���t:&Q�@������?܃�_s�~�x������0%����ַ�t��X�2�%�l��4����k��W��U�N� �L��z9ξ�<�\F�{+��b���t��*f"�Z�q#�^����&gU�KV�@�)0����/EDb��tY�zzq��g�gd������˯x9.��b-�bk���5�Qd���ĕr�?��c���J���u�����fA�M��׽�-�؄����Q��R��3��+_�j�YP�5����qI�"��cHP�s�I��3��$�����;nA�<'9���4����,���3���λ�r����;�x���G�Y�I�J��Ug�b<ͶRYӓ��`���2��������]k�{�溮7��%�o��
g�q�qT��3ڪ�
�P��
KͶq����т�E��^�뚰+�%����c���lŹ��DU�������V�[Ϲ�h�魭�!q�p�c�f[W�l�����<��nS�'C��4J6� ,�i�c ӣ)[2l�YZ���s���#S֪�d��#MWSǮs��n�:�!S��[짫a^�4�r)�td�B�O��Hm����esߩ]E���>�LS�'ʵ�`L�[\�	��7����	}�̰L�[& 4ZO�m�66m�m�6�m�f��vO���l[�}���|a��g����ZN巹�i�;����{'���z�үĩ#|WSr�|�I(���/�_�MD�Òr�9�Q�<y��l!N��������P04��?��-'}0�%�B%�q�vr�����[F_���3�^�>��M*D{d'��ײ8��ja�ԉK�4_�a�X~������V�,ܫ|e\�Qh�r^������V�m�w�SA�Op}���c�f_��Z�Kl�3��=�\����}"�0���վ@�^+}��oA	36�vxYчr��DMT��3]�(�$"۽ќސ������y��y�oY�w��X��[v���<�l���>C�*�G��È���S��I-�%G�5�;����5�09#��ͶE�e�!`0%�Z�T�+Yч��N��DyGx���p�ِ?��]��JmR��OC� ��r:ʄ;��$0�������5��e����*O�����k���&�, 1��!MF*7)���	�p��	�������$�����iT����U-b2Bף����(V]*��2��[R�־�SFC�~$%!��頳�|!�3�O#��p2 �j�ѭ�\N�� �`ݭ��K�x���������A�>FT獍g��4h�)�ߜ1�Ֆ֑=��g}�1�yw�k/�}"G�%-d��T�B0�j���
a���3��s��Z!8.؁�z�_<4�/��ȧ9?9�l�?�;e���*֖�����\B'��{�վjVa�$����L�To�oJM��@.�D�u�k�s������J|�@����KI��*ވS6ט�N�
o(U��VؠT7>.�BF}��'\��[J�<3�,�
�MO�i�f#~���M<���E�ǤeL���;T�Z"��&�hx.�t���eN�@���������#˜�j��Ϛ�.G������YQ@�cv
��!���t�B�97�	׊&�i��aՋ�oTXD�y%xi:؁�����8���}W����P�גF}p�HL��QRp�l=ϊ*ܺ~F���x��?��x��?jB�P���ٓf��!���8��WT�Z����bP6�=�1 +��<�u;R!gV=�>!�����*3��ztp��鵽[��\uJ�Q�r)��TE�Xa�F�0��%B��t>H^�,�m#�S��	2,k8���( �O�~x_r��8�/H������O��/X�>���>�0j�(`�I����p������,0��ˢz�5u�h���j���<`�TG�8�/�^5�^���h����y�UCl������u���5��O]N;�6�}�fҌٵSv�a�K�ĚY�ȶ�����#��O��8E�޷�ws���֓w��Lҋ���jBg�̽�<"N=:�]�гb�M�2��R���Os��yzCz�	����-�k�C�=�
J?tk�O ��xZѻw���3բؿ��u�i'ru�L8�M���A]z����n4Xu]�Ӟ�P4!�H5u͗	������)������\#a}�܇='�� �ߒ��{1o�vq�+Q�{#\�>Y�~���:��7l�:]$��!�}��� ж�)�R>.�a����g�s4O�q�����Vpc?��X����=Ro���(q�rH$�gi�xxl[$�"�&	z��ilJ�K̹����ǟ{�;�X�vڲ��`M�V�K�0L{~_�J��Mui47��*�o�ݳ6�* ����?<[{i�-K���3����l���B��g;2��A!d���I�w+�"n���V��܊S�H^��F.�\K8��6��
�܈u�h�[kUHYB�sS�����N�Gj<�z���'^��"�K!FM61��楅(6m�$U?Ʃ�'xbt�ʿ�ɵhN$>�?)l��U�Ԫ g.��9	 ip�^�hK��`c��M�L-�
�� �Iѐk*8W���,�S}9]}��,n��m`�O��dÁ��k�[�>���\��+�(�$Y�����v6�ȵz4:k*j��m���JmA�E���-a�u�o�Ai���P{��\��z��l�{��q��j���b�'vӑ O嬼g�4D�:|�ٟ�ū���]�\���h�^=/��6=>\�_���_�6���Pz��"���JJ�IO]�2�M1���}0��g���<K�	Ψ*A�{k�K>+�E5�w�O�
5���,qt��3aψ��u�=���͙b�H����,C�i�c��s�S���\�z�юe�=G���X�ΐ|)Fg���,J���F K G�ќ
���S�Ycd{C�	7>���ْ��/A����&N�9��ˎ*�f�����x���m=����Qui��.�����e�%�����̉�"��H�~~�0��?v>]-�̀���7��y ֓�5�CY��n�f��$��#0ƃ��N�y$_���V��L�O��_�96<`;ÎT[vR���c ���N�3�P��H@��[�&�{u=2.J�Nƶ�9��[	:��7�,�~�׋�l�2\�����,,���e�e��x����� � ��?��X�h��V��H���N��"�Ƿ\�<���3Y3���k�f���Џ}��[�e�M!"I�mt���^�4.d$��l��q�L��.��GGl���d�A欑=���%޿��U�W^>�v�=jD�y��lx�g��l&w<��0R�xrY�~6P�&݈�  �ö�rAR?q����槣�]��߃�PZ��������e)����"t�7�P��s�c����z�feo0�y��L����,�^'\�?F ��)uf���	����{�Pe�z{��ws�K�PL1��gY�cb%��\��>��	T�w%�7��Mqf���'��&t���x�/����O8���H����D�(렼@M�z�(�>�4��#�Э8��1��b���ܹM�B�����v�S�%F!Ȗ�H ����S��3�����5��tK~1~p�����1�qwf!Q�j����ong�6��}`���[����Q���쇠\���.�us�uD�g���q����#�@ȁ�FJ�8�͡�#+��d���B�|���`%����tkO�(c�	X9�+���ZJt�?����(��!�����y���\��`��b��}�î�'����+R 6�U1�PR�ZJ�Ů��r�aW�n(1���;�
W�����=[쉰�W�F�WL�����L�,����~"�:Y�H9�.܇i��c��N�O���.�m��&b��W80`�jR��
A L
1�
K&e�����N�>�1�`���~KM>G{����[�1��/C/.�^	LÂ�hM]�u-�����ґ%H�{ڲ��I���d�	�Ʈ�C�[5��(53V����x�KW0OmeyxY�M�"2y�Wo�yW����_$C�r����>�K��02q;�8�ZDf�Al����4P���D�V������b�4�e��pW��� �����_t��.ƱnJ�R _��ί��(�aBtEV�}���Y����~��D&V�<QS��|��>���g�.�&TS�a�\�����6��A��S2�ש�4^�8w��;r
D�I�[�n��%����l�F�C!��g�,��8�#&	U�>l�q�A8�vUu����֧q:깔�����m�7	1�nb]�TL�OR%�lؗo��<��i�
�[���"��(m�q8v�e������Z�ݒ�4y�x�SׇW�0��U���/�9�O��P
�aC�F��|@?�j���:KR�}�Lf���H�W���"�MP���n�������Kͫ�M�iY0�O�?/��n�rJ���,asbћ�8L����\2d��q��y��,�l<����(����g)p�v�$e�'亳�!I���z,�!��Kj/�,�A�0w�����A4�l��;0m����+�Q���~S\�Vg�-�O-E��ؖ�"V/?��a�fӣI�d!u\��(Fm�O���^�E����p%d9[n�O��B����T�ү���c'��L<�/o��~k�Q�����D�L�x�Ĵȱ��Y�H�	K+��џˋZ�SA�4_��\��*D�,BL���fV��Bc'�1�GD/|?-֬����6��M�ι��J�k�n^�&c�3gF(���1�#D�:�R��˪T����/_"�~6"�}"����MC�_%��FiN���%�J�o�]�>L<�0�Z4��:7�rĵ�O	�峈�H �9{���l�E�}ʕ�;8��c�&)����0%MVR0"�X���n�r;�&<OW1�g�&(Y9�ʍ�Ξ	��#��6�]�������<�k��r�l����nBs�u2������ؾԚ
�WY���7
F8�Z� �'�?�8mQ�o�L�����}M�k��+:B �ޟMd�ۍ�X���Jq;f�X�cm����g�K�i�Y��J����	����c$��b��k�x5.� I!�p����z�G���Yc��6?Mʓ�webdDm��s|��)���U����|���b�v>� �U��dƼ�"�E�~�RX!����WK�lDAx rk���.k5)���@h�<��c�;�m�o�
�1���\��ں�/{�]@�D���u�Ϗ鹁�6�v��jx�po�.���za?ے���֓?�1�� ;G,�by��eNB�Ӹ��0����d�v�s+A�fa��ã]8�C�)	�T��!m��pUwv�,�k.n�~�#
�N��c	?��?5�s׻�K�f��/C@ٰ�t�Lϖ��$���j��b����I+,f��y���3S����r������,���Q-����'�qѺ��A�w�C����;�v�m!,l�d���E=�x�3�&v��x�����S^�pݙׄ��x�["�ݍ�f͜��ƈre���Lr���@H�Ba�c Î2}ϭ�n�Y.�J�����[���	Q�\&_�r������ai���i�o��N��B��b^g�d�a��b)���D�fp����%��u zk4$�rY��z�j���/!ZfX��YAnڋ��|���w;(F�FV�B�j֒���Fp%��L���=u�=M�������7{C�Q8&�]ڛ;,5k���G�;�	��:���\Q�s�ocR�xٖÕj�=�N�2PBt�_Ĕ��^OkV*SǍ���|a������7���z��ak����s`�LF!��!���|��<%D���yJ��Hp�ȧ��� �tp�����⍿��<+e���E��V�R,�ɞf��X5*'{�8�����z��^�,����%����B�˪�G�c��׍v�|"�\*�,�,��(ϕ�]�^���v-����E~I���*�?΅�%��e�8Ń'˟�`��k;�+'%���lfz���y0��t�?���?/�i-
>��~���}��_Xb���u�*ܺZ@�=�T�X��Ȏ.�a�7�O#R��(F�{�GHʸ�od̯i�Ӎ����t���5���K�c��`���,�K(���x5yj�6������K���3�
�*�I瞜M��gG] �R��=��./`��B׶/D���9����x�Z�T�a'��X�&<����6Z���_���ZQ$�L��򗮮-:=����g1��1�#I���U{LL���_�hH͑h����ءJ;1|^�������dߠ�0{�^V�(�(V�V�������#�c�G��RG����CK7M�OyJHXJ����AN6�ZAv�CـJ�	|(^I��~0d��ð=T0�iL^�䭖���o��K1|c�XHaw9!o��I��9����?M��
�㏙"��h��
v���?�=���	��uV����le&d�Bt)Z&���񈧳L��4�?�ؙ����kk��,A�3�p���oP~x�S33��AMǇ����K�%�&C*�J��B�꠪�0h	Ї	5���l}|g��֗�&K��Qe�%��!
^N�`�����-j����k�Fl���s�>��#��L[~�x2W��8���a� F!�@�y��$�62Fc-�l�En�M}���T�,�a�xSL�s�	5�Pe���Q��1��w�r�ی�������$8��RC. ��"A���}��i�i��!�MN=��������9���6�4�w�~Y�F�L���=�jT��QU�w��Һ�,�8Z4���#�˘S%���T�f�}���;>��q'��/;�k~���8k���'�w������8�,%Y��UJ�9U�a0ud5����p�UvA��l=�0��>�UקW�p�f���*NpD��k�ᨚ� �������!$�Z!�ɗ$)��������~(oC�yUھO����;m|���o
��M�~'������S���`�)T[Ⱥ]�f��P�S
h(13>����Y��2�&�&s���.�ה�S0=����K�g���ઍ�G�|�I��^��x�,���I�6Ԡ��*3��9�����5�	Ϛƀ�$��Q뉺'���Z�
�(��EA��Xs����( �T(A�r�K�:����tpҢ�o�9Hh���g��n�G�&��n
�)-i
�T������ik��*(r��h��7ں�I���|��ן�R˱�����E<�}��)��<� "�Z.8vs�=�%���Km��	A�}�Vf,���5�`��6�,2��EѤ����?���9�����C��
7����3�
>�V��E["��T4�����x�N~�֗���`FQL�2#��وB�{�9����Y&@Q�7`miSڈ��f�^��As��71DDӵ�T���^g�V����5]�IƐ">8R�-�qU�[�c��l��U7��J"%\���䗋ּh�ģ,��K��7�����}ԙP`'��} >j|�il���|o��k/}��P��Z��g�����wBl�����/r�i֟7f]C}m��"�q��.@�[�|��b�
P X֛���<{����
�d���Ҭ�E��s?\���8wtc�����G�b�2��Wl���S�`=nz}L���-��Ǖ�4K��[�V�,�i�nz޸��-h���^d����nXV��i�֕[ST,����ߣg=⎛5���?�c���=l�A���z͖5P��P,gT�����E����Z���䤺�PM��_��&�ڵ���9ȑ!����K�YKp�\ޫn��M~CU���E�F0�ӽ{�f���Y\5kT��~[�N?�%(�{�a)�y�&Qc��Mʨ��IA��ϚDt(�T~V�Υ�?�E��7%�T�1x9�֕�d�(d��󮱨�����|�PS�~V�7�W
��.����$�s�aP��5#��������֨����7u���m�Ȉ��t�hݟ�?��ICEh�V�-�?�k�&+ wu&�8������r�����Ѽ�#�P]�D�y�-�&�Iƍ/�n^�>yB��B�#����W��8n4�~�{Ț⿦�9�_m2�_~nw��m}��|�
߆�b� 
�#fٝ���k�m?۽P���=Ȧ���^Gߵ���х\��d�w��g7�{�L��|��S��_$缲|=�v���wj���1������v{�w�#�	\WD=��'��S�
�a�娲)J^I��I����c�CZ��� ��H�.�$��Ӡ�hf�����n�V�B8���v�.�9Ƥ�Zvt��]k�÷o�s���&��&��[�e�lh�TC]aW k� K�8��zdz�O���@6V���?���jyq��������Pҕ�B���)��{T	��Ea��?��M��AAa��8��h�vXYA�M�&D�eBh�� �z,"p%����mTE2��_���k�Ӻ|_��Y�33����qT��[zw�ɤ���@r��X[�����)�B+O�����7^4��)X�\�Sى)�Քt:azm�������+�Y'�s����?{�
;�]
��,��-V(�z�v�
��U���\1��lԩ�n$��+��o�8f��n��)�b^sGk�����z����m�2�o��%�:-/�K��A8��;aY�ڌ$�C�U�ȼU�Ӹ��y��^?�`P֥�sF���6:K�)S�%��>�7&c��Z���)Ǖ��0������f�2��WQ
��`?�c&��TH��5)�݈�� ����Z	�̐���W����,.jE|B�[6�E"e�{��첰	]�:v^q6��5qI^pB�f�Z���a�Rr�v�0�țK/e���ћ��u�UAL�u,Xَr�=�
��
�i�^�,ǟ/������XF1~��Z�r�y��p��~{H<�΄�"�*�~��;�����F���I�XI�5��)�����Z��#�Hs���SN0-���r!_u��ɸ�8-�[ڇ�U-��Vzxv��1��oo>ƚ����s�a`��gK�V���s�xx�	+x�#�/aM����w���l�t��0�5�Y�v+���f̻�MLu���mme��+��6|F�QZu-+'R)���c֦[N����#-�=ӽ���9�4*��[N�O��ݬ�l$&~�.���n�^k�u%�Y,��+����'�-j�]6+��������L�K`��o.5MH��A�cڒ7DT0n���/��Ti'��$~��=����Y�����/����u6a�� ���@��%���cp�>�yvjiJ9��<��^��Jv\��k���~I��O�3t脮0�g�T��Z�r���{^��
<r�@}��r�۬����x_͐�}'an���y�Z�Gw����g����s����w�VP��~�2:o�|D��~f�|::�Q=�'9�Wa=N�.&�)�X�<��9��3�N,fR�3�*��B���(vv��ߩ4Ɉ(G."�x$[�?!����[&��zW $�C�t�E�3����}2�Hh��Rf؅X��A�Z�{+M���HI?$����t��Xܙ�k�N#\N��J�I���P��|�M���c��!!�9�Y�����j��ޫ{�je�ǻ��1=��X�<���7���,�ةШ~�b�Xk�LE���?}���1]U��g�RG�kjι��o�PŜ�x�x��q�����/����o�Q�k����ץ��+�XGcd�����8�;�����ط��K������Sw����4���d�eq��#��Z{
�gLɷ,�j�E�?���̪�H",�w[��a���h���������L<���U���������N�5*��~�!NH�G����L�����M�O:N��1��l�떒G�~��5a����3d!�{;��"��e��sKIK��X����eLez&2�����[�B��ٚ�V;S�8C�l�r}����9D���w}�7v�<����t�f�l(�mMʉ=�����=3�c�'��&�x߈+��IOsi��rR�ֹ�_6`�q����ӎ|U-�^�9`��P�s���`�2~g���>�|�����9��XO��J#��rK���E܉?��SZ�e���/ð"�V�������)q����1��*y�l���-��8�q��,1{r�C�u<	g��Hr/�^����+W���C��:+�nד��gT��dAz�$b�	��^��ϲL��g����:��ރ#>!�`��ș�Lب�8���W�x�0�P��N__��p� %��54�k���s�܉�uկ'�]n�4	��~�&�Ԗ�':-�nw��~h�Θ�@#����]��������p%̪�X�^�����_����D��:�e���u�+d�k����h"g{� ���.�D f��������|b��[2݁yry ����YG�y��d2�}n+�{HdS��#M1��V������G�n�0�T�2<%��Q��y����<���1k���cń�ă��aD��:��
�cu�����J�kv��@�,pʝk�]���|�O���J��:�}!�%i�gn����,�H��s�b�b	E;�B����.sEh ����C��0�]a�<a��%�.,�̋�a���f�K��v��C�?�B3%�_�`
�c5�.���G@��U;���_�+,����`��(�%�z�/t�W��,�D�;ֵ� 5&�ŒA@�p�kL�5�՞3T�6m0��RZ�k������w��,�fNZ�h�G�# U�W+t���v��2�+�T�s�,dyS&�߲I'[X�}�=z}܎y e�6m�G�������n�^h0X�p!��و���U��h���5�`SWh�N*�B��t�-ϸ�%I��.����72�<A��:��vYY�H���Mς��1��D����Jr%�}{w�Е W8�Q�W$�P��(�M�
��ˀ���gOB���?�����^Q��`^��/��}�E�����y��)���{U��ߨ�~n&k�H%D�&gl�aqj�I�%vkr�����|,$�<�<f�,i�:�*�����>���IU�!�jE�Y~���}�L��q�Q��pweM*��O�mG�OR��,���#�^K� y'��P�����?�sݹ�tƩ]����/}��"�m����KK���[�<lQ�xd�	(���~�$7���*��ۅ�_�;�2c�o=��B^�:�d���C(��Q��$�$��^�0�eI�J?fh�\{�_C�؀�Y�(���A:�³s����b9cB�H�B@�������@mʒ�(���<���Kɨ������b�3�
Re;��@�`@@�&�%"��c���������H��^S�V�|A�7̲RN��ڝ�>��AK�D�.�*��<�l`�|F!_Z��&op���I�۝(�	�Ǫ98��fRM��U�1W-K�X�s��{�H�'{��G.ŵ����9<6a�L�k�͜4Q�b�X�M����3����t
kƃ�p��v��xl52rl:R�C�ە����`���d���I�����z�nǆ
G�|��(�i�K��ڪ����I��`���^��{���M[��WuD��0'�~48~�  ���N�"�����ɶsm�����g�����<���	��W.*.�r涇��RMv:I\z��ր�Ir�-��v�LV��d��������Ǝ8�f�^��[C���d�(nC�W��@μn#��ۣ��&�����/�O8?��V��޻qdN}�z?8��`��`g�x��hTZ���5y�t@���
�Ky0j��?�:��6�!.��+rK�u;���y�̼K���n���uK�R�-�jrq�{U?CE�C%�����|��m=��l����S��G�i9|��
����I�����(^��Os� a0�M�g�.9K�G2g�@o`5�>-~>���ϵ�$Vkm�w���<>B�z� fT���N�іa���B�b+2���->���`� ۅo�p?t��>�1Y�%k_��_����L�=T�7����CO� ����;/mׅ�cn��st)F��3]G��w�N��A^�����&�ۙ{�����H7�-H�3Td"��S��$���͉����kMX��v`W�~ �Ju�K��zc���G��;W\M@Kpbo~��<�����l�uع�Ǳ?��A�
���W�C�>�,5��`z$��1��Fn\_{�����p9�]�k
9��+}QFo�򱳤�UC8b��;VWr=��"xR�!���Ǟ�Cy<;Qk���fJ6O��ը�������qdb=�t���$\��H�Z{N��}܃��s������a`�]�LԦ�x�����]�����P�˚{%ƈ+%
-�2����]a�YK�bb��8?"�$�Yk�u���㇐��J�R3��$�d��׿�G�eh�x/������|Ҵ�r�����H�b�͍�ޓ�]�������t"�b2�U1L(�����	,��b��[p��V�z%J�ÿ��n�P�QU'�e�$��7��	a�Q$?+�F�m���|�+�}ה�¡8��%�1g&�+�����*3�mr��y���G���UuF"�N���ձܒ:)jl7%h8э0}�~����#ak�h�њ�߈��@ekw�R�E��g�:/��CFUO�������"��bm�����׉�5��`��ς�}�S��8�q�׆
?h5'`x��i4;6�>spk������ ؉�6"��E1�:4�W����u��2.-��(�~��lj^HRR�l����� ��$[��P��)���c	�h�b?�	i�ek����t��R^5��\��(�4'��)h��gE�Z>���F؛K�m�X))&qI���������W���P��+d~�e��#A݃bSÞ`TPI��{L��+��;ϟ���[h&�&��h��z��%_֛D���F�.��$��S�@�s���Q�V������p�ϔ�8"�Dhl����&��&y�z����V�?�`7R���.�a�-1�RA�$�.@�� I�s��4W�Ҿ�; тC7|����]�/���a���a�E�����~�E )�X�S��܊ӏA�f���S
^/k �J�Z�����+9rd���Z�Ձ���vqv!�]DQ��-�knI��s�Qsu�]�|����� ���vy�@�)��ߝ���R�fl\��j�L��q u�����}�F@����y�j#�I͗Rݪ��J�0%Zjq�cc���3N����b-��Ё=�;�U����w[�S�r��ee����珐�Ą)�:}�����������<�7�]Ukmm<ʰ�Z���È��-m�Y�K�ꤻ��n�́��S�	����kRB��Q�In�����I�����)Z["��C믫H7ʰ,�@���٫~'�ן�����,�p������"�$Y���jÜ�\� ��#�JK�+6��!WLQ����?:
��|o��Ơ2~l�%ÄK~w�_ l�2l.�_ ��V����۳�]�+�} k���*�����-������[��d��%S!�H�+�Ӧ`D�[��+:�e��M-�pD�=I����(��촩k�Bz���)�`w �ԛ�r>q�b� �Ї|��[�~�_�o�4�W�~n�M� �"&�� �[�r�LBA9�ƒ�SYY�ؼ��5����oyB�D��m�D$��%���Q0���ũ���\�D��^R~ݍ����=���m۸��IVv->.�W��O�$���c	x23�&�4�ɫK���5�Z���tK��z�Gr�ͺ���� ���a�� ��(��^�M�Db��Ą8J�G��dY��HC�ș7D���P�Duy
�Q�aR���
yau�����KEߕ���4Wb-��n�]n��5c���J�O�|D�@���X�}���|�(���.G+3��
RVn#`��f��L��/9C�:�x�7V�f8! �*S��f
^d��ӑ�$C� X��.C���3x�ڐ��0�V�j����Q+{�;C%i_c&�2�,�el�B�;�{^�Sd��?��#Ο����<����6�u�W!:V_��^�6o�����9:���6���r������`�~d���shv�ߧ4	8B����h��o!�o��t�-����U��)������X�eh�t�#��	�69�/+m������C���RҦ��ɠ���Ѻ�{�xj�%����k�K�g�xS�ɸcl)T.3.�� %�Ԇ�B�UV�s�����S�Y,dx𦞎�1>>*�Ժ-B�$شxK�� gY�!��I(	(m(i�w.p-�	/�i�.s�9�r��VC&r�k:-���:�Zȏ��9�O�0�6�Do�a�ӆe�~�w����Q�?�RNM�w_ ���}� 6Ւ{�R��g)�)�B9u�,�=��.CI�|IA�a�39�AO���.ՎX�Rf��Op�4]��FpȍӀ_ۃ�����ى)� o[����_B�����VW�V������f^2����SЗ�S��M4%	��=;.��AZL4M��&��2h�$t�:vB���7����QHU9,𢆲1p)�����eF89dj�\���p���]���-]��TUv�ԣ�_e!����~��}����i%0�a���߮c֬�9����g'��)x���zw&�m
~ ��y�;�x.�ˊM����R��?̖:9
�h��B\�1>>�d�2�HB6�L�}Uz4wv��r�iyP_"��ۍX^�8�A�'�a�Q��7�5ߎ_A��u{n �����/U�~�,�k�R���9P�{�U�@��Ⴣ3U��;:�j}兒�騞������#���e`m[����gڗ��] 6$��0:�"����|P5�}s�cT�4��=�q���ٽ��Bn������[t\H��_�Ğ�1��=u������ �l&ɢ�w���v!�����t0k��j[�I�W=��&<؟�����C艼�؄p��F�pҨ��A�
�-�X�Vtmtc�q4���⒀<��)J��� �*�U���ډԉ��8]J�LE��2�f]z��������������"��� >��"�"E#��"]:firpж
Ǟ/�b����/��{�88�nK���3�b1X�@�WY߶	}���C�$���LԂ���ΐJGޤ��ҥ���9����1�Z�bj�>��.)+(�C�ܾU]�B��YӧTuQ��]	Y}�MѨ��Ys�>oX�߅>��3��mz�V ��PB�HDG�*V5��D���&�|�%�G�|;|L����W�Ax�/���Vx�Rvr��P/���o�BՌ��2���S-U�V�����I�o��K��$�ml�	Y��>�EmG��� 6RJ?\M��}R�D�x=�Z�h�d��xl���J��#yh�7��~4��K��SD��Pٞ�*���U�:n ������^;��d��4������e�:��v\c�8PZ���_[���z��{| ��H�}�]���-f����4��J��1�U}�Z+����:J��u��,���/���������i���r����|l�kͭ����-VS�����2q�)N^$�fm�����s�NM�P���[�HE�zY��V1|8�%�.{���k�ce)�{"��t���WjK�bU�=Y�@ԴS_��9�oP���9د4�!�R�?#E8&̾i�0ܴ���{ͽ�P�jTdPn�кG�E�!�/��g5����v��L`�>Fb~ö[���铽s9����:z�!���;�b<g#I����;��fg��-�5�R�uY�O���AJA'��æ�q&vVo�@�}]�ٺCj�<��_(�t�N�����Y:}�����[Uek��J+��Y��e�����^_0��4�i
"z���v)6T�y���""�`�t�՚2$uʲ͑Bp�:Vuğ�O�M��<���*�=@�
�%�: i��\K/R�'�
9��Ewo����kC��t��eH���ʢ�:���CՌ�m��By����g�M.��9�P�#��82�xaԴ=�}y��^V���~Gz-�|Jo�_�3z�� �H��y �Ζ����"��2�T$$h�1��ᆫ;#n�)��P.k@��3����n)<;h4�Z�d���>򐷢����x��7�<�hn8����(�*��J�\�'6$�4�>�3�.��Y���T)������M���S{���i'x�B0io� ����v�T|��hM[Y '��UN�f[{���"Y���V�S��h��  �mK��� k=��(;g���}��z��q��j��y6�G�fNE��,�k��)�52�.�`)��rn�2�=QfD^� ��.c(�� #���x�}���8;��I����H�Q�MS�K�@d4z5�	r4L7�m|�_�K�^Ȭ6�c�BW2w�K�^�����rC�Ovw�a�v��E=�0S��u}�U�R0�M���_#F�H���2�[@J�xKA���z^G<	�i���c��/Ch!�p1%��7V�Ƒ��6�]�����<w��v�+ yc��hAޖ�M���il�@o-"kr�<UK������OD��;��w<��]r&�I�G���2�桖w2ƍ�>7%k�~�q�]�Q����~AhEK�� y��^$C���{Md��Q�G����0�ĉ��7�<�zmNsWj�->>~�O�
q?6>::�,^v�҆��a�+��`�l��Ƃ�K���$�[���IpwHpw�k�5����?sgw_�|u��TG��z��$}����f��w���[u�T�����������=����p��H��S_i.IE����q>�e������g�#��o50�^�t8��l�Ź�mFuH�:�>B�� h3K#n�0���Y�݆կ�ynf��I�Wc��6:s[�#��QL��Q�8���'M�z��8+�����h:��b	���N�俗/s������	����_чX��F$�a�3X�hy&9��������`�r�Ҏ�+h(�g�d����G�@��1�ݲ�;�|�c�l�g�E����E�1*�T�B=̒�ᧃ�IXQ���>V�y�I3�����Dq`�����J�>}�>z�|l�o^�
�7ؚ�g��z�pZ���e0R<���(�����AN.�|��|����̒��J(ǳ!HN"�|({���e����5a����V�C�_+��"�⇔7�[�����2��*mL��7�i�^����"9T��-&`Y(1A?�?�"ԫ��1f���X�	�lT�l�ҹ��:����k�����9�0�?��Ij
��!F��0�N�� ���!/�N���䛦�f̞�߱�\��x�ey���&op�g�!�	�d���[�ؕ�� l����b��Һ>�X�(S.�
�w������|��*��� pT���"�{&E|���`
���%���`L3�Fu~E:���=-��qEEK?Ce�kDɷuX��lS��[��D_��c�g�cI�|��"�VZ%�a�����>��Z�i-ja�}ֽA��fu]?y�˴��r���eJ�-�m�Н��Z�C58Ec��ն�*kn��ka"���BWv�c����:��y]��3�E,J��ͷ��~o�T	��ۨKf�n4V&�q���kS��#U�n@��֫���U�<���8�j5�Y���t���*��6��X#��T_����5����,ߔ%F`}:�d�?�.!C��;����G
+n �G��T("�x�Ȏ�Sy��f�����o���Ⱦ|_vſ�_���K�wm��݀�uc#>�p�~��<|j���Sg����B����>�0��&�������#�OSlB����$-ny��YG0Lobu?�뮡��%Zɬ� &�?�(��p&MڴK~�����\5�:g� -�;�X��p$��+R�sGE����ļ|��t�9x?[H!K��eO����9<��L���B��:�<&|�SmbѾ?��TK]���)
[�|$s8FP0#R�1J���h�lSt��1e��fp�+	�c9T揗�j�`��&`�	D����w��
����!�,��� �;��U�o��iZ4�Ұ�����~�M�y��k��-��@�Z�l������"�6���}9op �0��I�?T���iR���QΖI>
�$9�Z��RXa§�o��0e��2',Ae��7+��Wk����J�J%�тnÞ`�I��༑�H1ǻ!�i̿X� (�/�zS�/��'4�!6�LvX�B(��xBid�m?8�-�8fY䭎y@����o�������a���f�$����ν�or�c֬\Q�+�)eux�[�H��y�������x�̓+vm� 4����=1��b��D>�:hT>�nw_�C#�B?�-X�&�.�=f ��q�����-�2�+�m�KY�H]C���V<���*�ؾ�H�(130��<�W�h���ש�JU��2���<��l5��[Ϲ��'��]���a�zO^�
��(����Ν�����x�d,l�$G�GD����YpݹEa���e��P�i5�S֐Y�^\¯YF_4X͕#!4g'�H��з���R�Ä#!!����se��C<�z}ɀ�ı���3��)Actyy�Ѻl����u[���$]8V��!%?�l,��C%?��k�?O�l�n�B;p*�fl�������BSN<����'�̆����ʬ�g(=��qhpQ�|�ɾ�MRP��A\���$R`l3�b[�ZL[7�?t����¯�.R��
�S��� T��-?�x�$��G5>�Iᡉ`1����:U�,͡���`��r��?ʭTSт�`y6�)֝���1���u\`1UoX-Z��g�}��QT���)���Ӄ����x�i#Sa@�Ai̐R��_)�e3^���T팴��%Lj<�r��4�FХCz�a=0���I�7H��f���s�!i>�~(��n�x��`�?]�0�2�7O_��%� q�a�	^�faK�)���Jj�2��+ވ�x��_��$"�{2�;�WuP9�[��+Gt���ή�VJ��K�̮)Q_���
H.k@�EG2�Y���GN�ҿ������m�>�j'AD}
�E1�\j4��`�]�h�7����Em�N���
���D	��� ���۸2�����開T֏��L�ڛ��Y���TL���2/�'P�_���E��I��Iʘ�땋�z�Hk�I�#N�&B�H�IN�p��̎X�ÿ��m."`��9޶Ԩ�fK�}����ւ�����^�-�����9��%��Dr=���&rRΛ��ƪC��ec��1�`���OQ�2�c��ʘ.�"�Dd� ��=�g��ӄ.�H�rp�5�툆<W �b��e�����"����2;~����:�ET�<�.%}�#EQC�-�+����˛i����f����f����`p����W�w�}�^��!n�)ԗL�d>�A�fd8d�ݚ���B�˕��ڀ-*>��v����+���J�d�����ɏ���v�?m�[���LhB�cgRo��-~?��>+?" �jNtL,��^_�ϧ��8�F�:�hQ[�^79As��
�s*�����Y���d�q��.�ȿ3iL�l5�]�ڣ�WD�di�e��[B�9N;�Gȹ�Rbמ�g�� � %�\��;��uY���̵�2�EY}�μW!��k�+Y0Vy@���`?
�lݏ��u��X�� �ּ����-=��*�m�����%-!��m0�b$�� �8R��f�?
�&>�9�Žb��"�<�1�*�����7�9���:�����+��#"�u/��j�|6ȥ)(�'�<� ;�+7�8�p����~;��$FV)�"�
.7��V�h|M�ԗU���qdk��3ߖH18!�6��%�=�T_�Y��v>���ϔJ�m��`5[���L�,+���ֿ��}5��`<�?�0��0�FQ3~��H�Ɣ�AR�fP���(���6M]f�C\���#��ZF��E.�P<l�J*���S�'�P�!�Q �F�A��� ����,.�klbݫY��*t@0�f�����h2��`&�b3(}����^w)��jx�:�SG����uY8�aco<����S:e
��0����ł7p�5k�"��oj���?���8m�p���	��c�|��C}a5t���S�wy�l��� t7�����r�p�7�Y�v�T7�����D�IG��������r����u�����9w���owfL����=��U��A��s�A�%���m�8�����,��ANJ���|k���Q�("IIX$l���'@�!����i`��N�ھ+՟p�y%\t��ϲ9�x�J/�n�y�Y���J���k?D�Nc헭����hc�v6�c(�ϒ��[{"�[�׎hխi١2=��b&-�ݐJ�$���v��bG\N���)�֜-`9���-�սֳ��HS���ܠm��Jy�F�2m�������n5q%R�_�?��O:@>���h<����ޟ���p�2Do��eV�8m��hպE��ˈ�dn���o���N(0}��b�����YQg	@䠿70��i�]rm@��B8�o]�l��߶���A(�!:?�e���ܙ>��B��~�g2�=�o�����qS�4ws�ig#������\��/x1C'��d��7�[��������U:9�	���G���,�
ѵκ��c����^�L����=�A7E������A��k�2�9(�m�S�4���@�?�����n�^�y��+̡<�+y�;�����-���)�h�n7���V���4��?1:���r:�1)|1y*|Ѯ�%�f��� �F�T��:��eiMLbz�Teꃖ�}����í*�O2YN�ʓ��w�B�K�j��8���.��J0ፉ�P��?*r+�x�9������(-6/��e�SD8�+����t?�yJF�/Z�諻c��k�������y�<̀�&��|>�9A���4n�����#�����
/�ZB2ig+v*E<��_�$S°������� y�FIh!�~�c;���N�b9m&R]W�����?|�ג��s�SK��o�XenOF�r�if����d���QR�����q�W�����g�9��zy���%�ikh�88�D&"f�t�@u!UQ���\b�N�~1�!*p����c�����wO,`�g�����9�)����ʈ2�+�pKp}J��/����@�G�p�v�����@8X>�x⍛�V����<Ux��/>��}���Ax�:0��yR��ş�а՝J�ʿ!�~~�Z4r�
x8�l��h�g�i��<�2	��!r[މ����T+=�7��w&�����Q�3֫�g䖵�|}�^�[��r����z)��pr� 9� ���J�<�����V�-�y!��=ھd\�h��&�EA���T���l�-�8q�M���ϯ Y�n"�)��ݮ�[� T��~�߮c�~;#�d��+�"%�X���'��3�6m-�c 3�����u�j��
:��O���)�`�L�yI7I�U���g&���F��ݥ>�7$�Q���g�5N�y$����q�H�����;������1�Wz����a6�v`3rQ^�(}v4)~i�f��[���_4�"k�Mv��B����\k/,��@�n]���$�%��?�=�y�ϩ�s\`4�h�VSJ3�N�ķ�n�~�t�7�v�]qPD���[�>��Db<�c|H?��b����)A�
.�l�A�&��Ty/qI6���eN�G��oԘ��-������@�l����l��#ʮ�/sa�����2�G@SSb.X��6�ֲ���72R�&�M|8�?�gR����L�L��;��`�L�ލ9�vN40�A��>¶!�������5��K��Ǯ~Br{��vGk��)v���H9�X+��λj��G��ͺ��ȠO����T9^S��i����{@#�{j�o�>J8+_����5>��*�(�y�du����gQ%�ob������U0M�I��!�p���v
�e:R��|�H�I`�#�7��}����t���z�ŋ쀞"�yAÄ��Y�J����3�Q=�l6%_΄7%�mPEE��{�ǋ$�Nh� ��p���(�"%pv�v�*%)�NX�U�?�G ��%�Ҽ���At��P~�I��L_̋��|k��NEZa���%�KC��p*�+�h�|-�'�c�{@�ȵ{d5��m'�����鋀��8�w��e7����  �e��иQJ��+63�H��h �9��`GU9ƒNbg!a���&奨$���K��S#��OR���)�W��u�%:H�NQڊ�K�([�����\��F���������ћn��C�\#G��֒}RD��ZW����Wi�ԓ�f�3z2�*tR#kt��G��u#����F��bM����+J��m,���D�IY4�>�.��'���hN�1��X5ˆV�d�Z���J@'b*X�8��K��9�#��⏳I�^��:)�
��,��_�6��lY�ߵcP*��N�V�wj$��Y�����O���I�!�����}.�c�(r� �Z�j�D;e�D|'Vq8��BT���/�	v� �o���G��O<;6�aU��~�S���:�G[D�Dc�z�D�D�s<&��0Q_������İ?#�Oh�l���7H�JsY��S��YΔ3�.���kD9pYۺ��܌b�8+EZ��ԡ��9%e�ꙗ|�q�Yd%�#��,'�V��Ø��:�V�"�x!|*�	"��k�%�by9b�7 F�2�ā_�'�:=x��S�r�����|�1JxC�p�[�X
��+o�A�2Q������|�U�Ej�yE���$��Լ���%�xF��Z�d�_8Q0���_{�� K��[����S��A���D�����,��2ߥ�?���<#����"���we�U.�_�G��3�|C��c�c�^k�X��N~��uh���aC�m� Ϻ�^J�>�%��擢ּ���1*߿#~�/ϧ#��d3��Ny�~� ��D"�yEO.���U?*�y��4q�ۜ/GU~>���mR�����F�:QW�=aҬ4�3(&L���'�ೠ�;j��ec���LJ��DpAJ���(�GiFa";ƃM�b�>k�����ǠF7�#���θW�9-_�m8��2���h`�G�%������;>���;���'���,�����FZ�B~�A�M�P}�l�hV0��%��:���&�E���+���V��Udq�p���)���iL���ה�2��a�8J~(��Q���Q��jb?2Z�>�T|�ܬ�ʭ�K�`g(1��Y(�O!i����������A���/~xl��}qsm �"|&l��&�+�S�e=~��<ZVp={�����
�ˊO�6�v{�m�f�
>	�CZ�D)u�|�I���u�[����U��*�����6�u�P�b�Y�qyjQ�!WJKr���T�:]WL�P�b�u*��0��ԏP|�B���V���5l��CQG���M#En8\�K�<���r[s`]}�-��Tf埊��x����#+LI��v��v������f4����ݏ~_�TG�kmW
��ǹ�#\X��!UvQ]�Hh�}A�}}�a�,u��ߴ�J�t��X2�[1��Gg�'�(�+��O�^c��0���E���\m�8�/���j�� 	�gvZS��eȺG-���~�Wv� {o-(-
�iq�d�eo$e��WT)UH��Q\�~&��
_��b��
�c:�dq��4	�X
�[��ШY�GU�DL9F�7c?@�H��:0Z��e�`���+;Qo}�O���Z�̜!��/�ܷ�*�r����iK)pB���@Y��2K@��.v���ȩ���t��Q��z���Q4���'����q���M���k�>��ѯ�-�z�z�!�ON=����G�j�!	�,i���;�1��J�Ό���@=(d�H��0�#?�C�Q���
@��9L�|qx �@���Ujc�0�V����c��p�����0���3�A��b#���2ѓ	C��'�T���o���j���(A5�߇�i��D z*c�Y(SN���7�4��v}��6i��?��P�}۩6�V-cK����/���cS��}s��,�P��s:�c���P
��p���)O��5�OE/L*_�h\^��8�*�����"�GG�nk,�"����uxB�+G@����ڛn�Z�Y�oF�E#Vb7jY%`�f��glv�z�?m*c��>��{�����y?�X>#�E�tD���%�� �,X\	��)������|����s}���5��L��hn��������.r�Щ�Fi�%�]��
�9��)���{�����7{<|V���/��S�X3�Z����xP\�����LF�x|�/�h��v�r��q�wV��� �|C�
-<-J���H[CZ��
AjQ[HsH�ia9@-��M?�:Ӣ��8t�]��NE�Ю��-:�Rn�k��B������D�� _b��r��U���{�ٖ�?��VG
l��V�t ���ĭ �-����͹���=޾�Ҿ)� s8Q��L��o��}��1Gp���}�gp�b!K�8jƑg��us�^;����{$^��:��/B��A�(��qy���UY|S=ۼEᣳ��*���f�\�ٮx<��*2�)��#�!�V���v,���bLU�����li��V��Ō#q��
e��T��{S� ��&/x�1O������	%����}4�])���v�����гr��U����3��׃ԋ�7����$a�Ol;������p��o�׮Vz�G��!i��j��z�CQm�>��w~�]F�}�%��(���["� �c
����h�N����0n;�����GJ�=����`�B���C�;NGGG�i�ʲ�x�E��Fj�o-Ĩ�R�=b]����������>��o���g�|0:�o��L�x�z��F<��48�\������x�o�e���`r����rn}�������g�m,���D樝4߄Ɗ_��.��u$�//�b�;�5�O8zXBG��_�8Z_x�n��=.?dN���;U�Ê=��Z8Z�X�	�1O	8vݢ�>?��NӴ^��n�d�;�=�>�~��Y���H(!!��ѝ�q�	1��Zݰ(yM����{��z�ڹ*�@�<� ՞�.��`Bbbb���x*�ӝ�`K��p�z�`��T�E�����;i`��t���W�2#$jᯧ�}�CI�B��GD����O��**p�k�U2d���!�A�r��/���q'$��o��OBQ�4�X:=U�~��,O�>g t3��d��Е���OZa�@SS<ɿM#���o5'��	��%1�%�a�d�g���:p�hB������7�l>��d�W}6�7�@0�K�&�Z�m�K�Ei�
�K���_| 4C��̼�(�E��D�;��[���7h/�BW�6�G���]{�fîV(�-��?���B)uh����`�T��s��u�?hO�:I��:�e4�&9��8o0b���V�\�
)��7U��ƈ�hXa�����%Ņq�> ��
qa����&ؒ}�����q������a��]O�z���?��ɍ�����9���1��Bu���\����#�y�����6�۱L�;4����ٍ69X�F"��L�u�G�����n�~��ܜQ��1��uj�F��G��!��?n`"�O�C���8>))y���=�|�ǯ�ՠ��"���������J�[w��?�|��ZFoYK��)�m�s�K�Ϣ{�b�e�)�^���D���ѫ�V��� |׌l}���$E�NU�תR��чJ��'���.,ņ~]G_�qyͮ���O=0w��q�ވ2����_2qedqB���"���h�2���Q���p�(�&�:��\_��T��d����p�q^�̩I;�ڨ�l�}�Ug�'Y��~�U�ؒ{���Ӵ��T���J,8#�c����T#��h?s����[/VI�����{f�֕s"��sc���k�3P�9��)A���b`����^��j���\�e��6)�n�X5����2y����ҕp�Gb���~-��)�<���}�'rh�qH\�!M�ҿ�D<�;�p����ކ�*i����ŏL*�}��Z��z� 1����9��O/�#!T�Q䁘�%�ci��]H��D�5؋���//Hmϲ|f�ٵ#���_��)F S�1��7�������|���r���^ �ft�g�HM~�>5�z�6��#|�5ñ�J�OMN7܍��;(��ZA�C�O�J� k������.�y�	�ڽ���#h�(���_���ezN�L�+���G[�8����z-�ڴ����~B��N��O➧�i����?&�d$���&�U
#h{���o�}4w[�Cƍ�s�'�8�ˀ/٣{��y�r���怵@�������S ��*_������N1"Lvk=Q����%����hP!po��aBy
�x�Ƽx{�ݒ~X!O��!�H����卑ýF��$���iM����j6M:1�-MP���c�Ԋ����av�f�iD5�@����t��f颪�N�x&a��
�u3 5~���rE���c]�ky�iF�(�S��ї�\�U���>j	�;�;���0#ٌ��T�8ղ��Ġ�?!�o_��u��&Y{����%k��\͖�'F/'�^���&�Wl��z]�t���(�d7�r��vY��0v�@`���lɊ*^�����圍�\�`����*�Ql��l�o�\Ɂ|B����̕��YZ���l��PO�XI�s���d+�E˙v���3���+f��K5���o	�g0H�^ �-�Lu.]�*\�������Y�惍�r@cBH��́�pL�d�e[��:�]F�����V�5�W��C]���p�E2�шC���Fn��������C��]GD�ڄ�����M�b#y5y$lz����e�|k����kۑ�i�ʁ���.:��P-a�@$��R����u�_[͏`�1b:��@nK���X)��a�M,28��[����b�/��Rﯶ_��Yh�Xǵ��:�}mt��R��m�d�辕H��d�d&�lQ�ϡ�<�*}�
��VE�c�E�Y��f�	�-�M�旉b��*eOr�?me���mjڪ�M�����7㨰�xnd/�i!���g��a�N�E�p�i��	�#�p�,D�H4���ԦN�X֎$�B��*]����h����=������\��JU�p���c,w�vz�
'�����)�$�~���P���f�4�v�b�S�E8�F��k�����y.��D�r�;y�;'*��vr��:L�c)����Y���0��A�]N�O���l�7�|Z�]�^�J�|�^��u0#��o�]�bF��psP�4�����^�-�Y��,W�/�0�� ^��CbDX�J]n�dG}u�ޣ?�@�l|gh�	���ަW���ws�������Sh��0�㮍�4a��uH'E��
KM��=o��������
8�JV�w�+M�
?����Bo�/�`<_l)(χmV�����u�aa�J����>���K2�A����s�Ʋ���hT��[4��5��F�&̆,����_"Ｚl��ȻOEMkx��M��	v��ϋ�	���y�����Ue�L�/ު̋�k�-JeA��W,�~�]a�ʚ�aCI��%Ӎ)%�����V����qM�\�2�*�K�rm��h���pfY��n�x�g�Lڮ���_���*./7X:@����0=�II \�Pp��Go��U���B�_�&�Y�^��b���0'o��<02��*-I4%o���{_�~�l����y?U�V{��l�:6����!�^�kߪ,�q����V�[��V%Dć�ٹ}�C�v�l�� �b ~�l�ݒm}ˏ#P����F�S�{\��;0-w���

��n qZ�kqr
��t}+4�v$��I[�伕"���
��KZ����U��$�+M��D��c��İP���֗3�	���qZoGX[�ig�KO�++B��h �B�����f!'<�>��#� \1�b}�SE�a	���&eq����~���:�JI�&���ldNd��	��e_ݦ�R��J��<�+�����w�����$z�{-�ܟZ�nes������E�g��jT#����w�wN$,��;?��s�%��xFh綇Jw��B�Q�4g��ʙ�J�0~,0�\F�X�8�F���s���~��&Ɉ�6���:���g��.qEY��H/�~ɽ��_��B�8[�nR2�}T��lـ/�o�"="�`�9�����ܲC���)U���d��\ѷe��i�IT.�ϜR,Rn������=��D�)N�Dh���Rņ�0Z�X�����Tc� a�iЊ�	WQa1U"kH�;ϧ�/8p."�F/���h`:�r��H����H��#��c3�����ϗd�>H���c�>Q�:Q�B�Q�_`���=���<<@�r��Y�q�~j��au>X�9��1���~��]���pS7{4Yp�zY<�z�ǃ�n���o�	+%!�(�H7B2TSFB��1���A�_�v��(�]�p���`��z8~$F��I:��Gӂ�:�O�R�B�1��Ge�3qrT�b- II}L�:�T0�{gD�R���`�%�g�^<�@��5���p��㟯���p�r9J�+~�`w�f��8]m��S{ �'�����n���p�����a���ͣ��R�5����� F���P��O#�}}/�9k4]ҮK
,�Q$%}�/�����c"�׳�p�3�����qS�ǋ�1��N��q�PN҈хm�&�u�֚Dp���3�*��l�-;�-�yԴ�4�`aYo�����6��p���sJE�gMr���?���5˵�@�hH�/FK��ٹ`:�\F�����B*�F9.Xݼ{RQ�t�|Iݙ-l2J�N�W!]��;,��̡�Hu�C��Ԉ,{��ft�g=������c��x��^�\���j{K��6�0�u�Osm,F��nO�:C����_F��uq����:XӪ��*33R���g���
E��	���;p��a�qcvښ�n~M���;\��~-���0<o���^�g������¹���C��������!�Q��E7�����aΖ���6��`��ʺ�˥�G6X��̣��0{�>cT��B>5��4
�%cۖ���=��C�;�o޴M�_E��c����RΖ0���#���>����/������u'i���^a3(I]RETb+z�ʋGԸM[�#�Xഝo!�Τ~J�#�r�$��|W�Y�43D�c@t1���W3?T:m��R���J�;Բ����w�`_�3�%E�{��a{����%�z������^`@@j=��m�q����6�g�B��k�d�	����=ȁ��4�͝��i%�j\g�����y��U�$1����jqs�Y'�=��m����H�I�����{�ٟg�|�]W����;�F�g��� ��z�5��NF�UC�t��2	�e\�k���i��y�	���Ӗ3׸o��v��/�SHS��^m�m��G`�61�.ҡS#��M���|���c¹�{!�������1��A���I1t���Q��}���_��@�@���jG�:��yL4ҷq�#�xVu��t�[h��4���m�l��&,�_V�Ǎp��?�f�0A��(E�&u,wN��:=oy�{̰nd|��%�b�o �UB�:�����]�z�o>��`$���z������j�k{E=Ů�CʂI[,���bl��ŵ٪���՘�锨ܑz��*�6���ՠv��D��̲ �A�
6��`��7ſ�Z-���R���fݘи\+��#�;W��(-X7�C#>	��5�B�,:�Y������n@6Td��o����c��:�}teϜ\�-��U��������v�Fk�*������I�1D�X��a�E��8�C|W;Q�#?�TkB�TEF(��+ʔ�t���XO��j��[H�^�0L�\�`�me+�|{�0�?���c�PdzӀ8����Ӣ��pp^+�S ��e�Z  Q�R9��{\�	��n�4��/K=��`t
�MJ}=m�J�� {z*�4:ΐU�lh��/vL�i����{�UFO��n���n����j����%�b���2h���S����H~p0'����A'�y&��������p}��<l��z2�w1q�U����m�k���l8F���ՠ�F3D}8���v=��]~�xq3���]~��k����^���Ъ�U���
�r�6���u.�{�ڧǦ�m����q�Q	�$��R����N���[XLC�7�ߤE�پ棢��D#5����4�#u��V�x��)ҧ���]��[����XF]�VC��;�o�'��a�*�������=oVf�<_���\׆���0�8�К&�� �K1�����5�}�OS�q���[ض�)��xhD�{eff��;��8���Ь�E𿛱,h3w_bΘk��H��� �48L`�>}6�#�,+�(��6��ʅ�vB�H�3v�Do@���T�x�jv<EP�iS�^}|h��N�Hh����G�
v�Y2���
��Cz�9�_���V�vI({�v��`�2��Y��K� ���}}Ԋҹ<wձ�{s����RsF#L���@,���<�B�����@�=��#�L�"��`��2��3N�La%\��� �d�:�VӋQ��6!�G!�mm��f'Ċ�GT�+U�ܼ�HX��ñ��Ϻ
*�B8ۥ툒<X��Zv�h(���5���x)u�a�6�����H�����i�-ue((��ܲ`rb�q���`��L�����l���U�_B��Ea]AQ?������XʱU�}���0�Va��a����]�e5��u��D>��>���e�g'�?-*z�?m�O�2���D`(���7���M�!j�*���: _�T�ʮI2C�K����\kh�kWD�Iq�(��`t}DO4
�4a6��;vE���8��H�\�H<�C��B�7�N���,7L"��+*��k�U	?����#�r��R��%	��L�k�^oЗ�I��A.���=7q+�@5���?!z�����~o�M����{�EL���W�-a����E87C�=Q�S
$$v��]��fE��̔�֛��3=B�����Y���p��: ��ЉC�'����2�Ь���8��Q�z3+�ذ���zI`B
�y�P�kӽ��xm�Ѩv�4�QOU�[�9�3���1_+����
��Xz?.�!�$ ����<���5���������
�|�DCۙdn�Cd����582J��sq��'�ܘHI��&V4L)�:^�l|V����_�S���$zg\7���?�B���35�,�����B�Ӂ[�,/F��v,u�)�p��q��S�pe��m��q����t7��"]76��g�QE{�X	ҩ	`���:NM�" $"{�b_/�bfV���I��:�KHۨ/�����iy��vI~d��*#p��Ō��П��$]�ݤ����Ӊ���<�w�����p0;.�qI4�^a/?��K��}���j(�&'&�L�7!��SW��4ˡ���2LO�%�u��sZa������P�z����Z�ä.��Y�]M��4[CE���i�L���'��_���<�.7g���Ht����
т������,��o26�h���T�Pix�0#>��}j�%�	�F��!���Ϙp�`D���=u5��hg <O/.f�_X>�~?����d�U��*�\8��0<�rs � "q����k�?utX�,� ގ��-�����r��A�Μ��`#��QÞ��O/g<���������-�S�3��A���ߒ3�`Ng��e��C'���te��P�T�7�/+�����k:2�D��x�IA@<o��'�G�H��"~�&c^���]A��r�L���iM:���7�'�`>T�m!9����X��������������Ȟ�΢��m�g���%�]R){�@�>����˹3���8�>E�<�N��þ�����L����X�U�~�y�ͬe!��Se���XF�}ɮ�pF@J��ٯI�M��BQ�@�T�
��ΐ&��uO�[̲�J�2��(�����Q�l����jAV2��%&]"u�N��ؚyr�qa1\��X���#�AZ�b�Y�$>�X��LH��dn�e�#�&挀#ɂѸ3�K{�K�u�9K�
��---oh�4���7?�l�� �,.-,�=%T�t���z�%~���������{L$�Ղdɱ�B
�P��j��
�׫��$|YǕ�[q$W�ĩ%
B-���КG0�~� Ksr�(w�y��w.S�-=���7��u*�X��m����-`X����[��k9:��Mw����Pd�G��$'���3d-�L�q:QYO��i~���Հ�"��E3mAv	�P������3>��5��[�����6��&�+��<�9���p ]�7+��l�IeŜ��o` ���� s� !�p�"2&Y�UV��2��P�ٝ[�X���X��!"HQ)qC.D2�����wB�.U��~����� �h :���@��M�x`�_ :�P��%�M��*���!hנ�#�������Nb���=��+R����T[P��4s.�$s�Q��ps.0�$$˷g4��ua�~�Z1r!���߭-��dPw�v��F`��p�`~�zF��/C���	˨Dd��t���p'��:&���֑��ޫ�����%��5�.��N���"Y��#�,���rl�8=Fy�Ъ��VoI�P�q��1q��9i��x�*c�:�?}.���i8����TAZ�D`�V?3� �Ve��&����T�G��i�lKk5w�O��;>�$�g6F�E�3��<}!V!������8����l]C!�p�����/4��w	�,@ᮅN� �;����޽/��s>�+c�n���84�A:
K���J.@y脻�o�{��L' ^~}�P��1OK���Ru���<#6?�z��e��c_Ő~"`�YNɯ�%�r�62j~/�Y�ޭ�+z������O���m�Lx��ٯ�A�B�6�+N��ڀ�����#B�e�)�]��ǯ�8p���˴5�֑r��{�<��?`�"�V��_���ݭ�k�$ǘV��{����z��D������X|Ǭ^%����*���ؿ��blJ���Y,�EY�AU7 ���݃�_@�Jl�jTÄ�\����۳ǾhB�u��!�����]#����,#$jƔ4�Ղ��ݪ��wg�pי$��sZ�qp3��g
q��0а��8TG���;��Q�d����1�odmDU��!m���1��T�?���_�Ѳ��%�)����u�����'l�'v� '��#�}��U���ٴ`�5n��<O �En�[�M&�6���c������n������#�*y��I��_`ߥ���f����V|ܠ,����#p\�۞E� f�jc@d�;�n��i1i����LB��<��@Ɣ�5���ؘ�l��
�R�<�uD]�����
�/Q?M�l�����3m���5����e7�E�h+ܦ�����ak�a�|�Wy����������P
^�{�;p�-tFH��A�$����b�4�/3��RX~g�=�T��+�A���O^��w����1h��q͞Ƞ�[�B��_��Jf��&���9C��X�.V;	���Я����i��hl�}vơ�^�����篫ꦯ9�����ϑAX'�X�7
�yr��5���� ��f�@b����ae��f��|X�_����8V(]���y�XT�T`�)-��Hz�3U�RM��f�B1�o��Q�ӡ�*���4��7˥��٣�e��H��@Ѥ��s���y���_�w�:�_A�9�"5��rj�����`�����3�|���΋9���~���_��|J�dҖ����1�B:z����\S�o�XF����A��4�Eyw���"���]J!���3?zg|�wh58���|hDޟ�n��x�9���v��Ʌ�6?���j��.W~�Z��Pq����yU�g^͓�^cX,ʰ ���M��|:���.(d_�qz L��,�<��'�GIkcl�H?*x=�<}�O+瓠Hܑ4�R��ءq�x�v��ҁ��ޗ���=�qG���$���[4*u��T�?M���D>@�՚��	�6����f���������yRM��Pr����9"�aNO� �]��}Lw�?��R�p.]>�z�*��$vΤ�HQ���cJ�2��Þ���\��*ʹ�
&f#|��;úђ���EN�F�󛻸��-`�s^�}w�t� ���;
y��"��)x������":&��Yi�H�e� h�[��2"�'
_��>��	vHɴ��еlO�]b׵pgjx��Q�������	
��p&=�=�g�T�/p�o�X?�b��łB�!r�Y\=���͋=X���[�
�R�y3�b?�l!��?��v�!#ⷊa��7^&N������l3���ʓd�l��O5�M�d&�C%�4����s9/_ݮ���=;�7r���񘑏H:4w���01�j��F��+N/B�����U��y⏪ɼ!�x�r*���3	�AH9dA�j���v��>�;��x���%a�h(�S/�r�_�
�$��)��O\k������ޠ��rXK��9I%��K�x�$�BzʠI����q�`��J�q�$�w�^m�uw�7���A����x	%*�S���L�K/�J��-F����Z$�������Z4ZW�L�}Qtw^b�����QP.���8�����c,Oaw0����<�����]�LyO�<��B�����rKlmUA�C����+����.D ����A��M�!����$�'iz�K����66+���fn��v���
�f?wA���Ԕ&���op��U9���W)�`v���fಶ˯c���>9ro�����J[���-Px�WLAّ/G�����V!vf���֌�`�.H,��!t�[��]�r�^��B+��.l�ޱP��6g�O�à�ՐF6��g������2i`�l�<h)71&5<���Vײ_�L��=án�8�C�6�J�N��47�;c���W��E??��k�Sjɬ�0=���4�L�x\;,yO,Ic�ܯ���;P%��{�|��Ǚ��|38��i�yv| �x�t�L��$N����6)lm]�X�6����sk{>�-t[`�P��[��Uc���zC�j�pq��LC��I����a��;�,��Z,��Mך��8h��<BFq#s��"T��~��.��˞n� �>:B��oN���T*��L�����\�"��:����/���"ą����r���a#�%~�J$lf��Fa��vjȝ--<L�a�60!��y�J�L��h3tw/���SE@7d)C�d�I���%��B��/���[wh0}�ã�l���JH�Z�A�r(�^��g^/����W[��8�S�0����gr�G���Ʉ#�e���Gq2�X��Ш����{��D��
�[ٿ>�Q��pA��m`�������C=5�,�Y��96$B�,��A�Q�v��_߸o�+r�y�XG���p�"�u��3���)��t�f:X�QZVz����_��|Hz��$�C��L[�؅��U)�)e�s� �H�m�n��uA�o�w��B�A��?ZWWy"��*�d����(���G@���+ln�˻��Z�8��M�(>g�r�qr���y�.[߿���]=��ݻ���v߯�׹��֜��6�j��1��$���KTm��3Qܺ�����X���]�ee�����=� �z��`�}Ӄ�x�EN^~�����Z<t�������J��tM;�K��w�nf������,Z����Q*2�F�X�Ŭ��XZ��:��A��kw����B����0�<'��Zk��p*[����3Q�v75L�3m]o5YR��Gjq?�Ő�o�G����!��pD�@+�̱O���\����� ї�p!T��T+U��	�2u��}�%o�~�B��G:�U���O���B�S��߇���33?[�kl�r=;g���؀�g%�$Q��k�&��%��}M�4f��\Bz0�C��_��-������aҬd,�
�$J-M����&N�-�ࡋ�GǪ�9\밤���h�bSHW�p��Q<�+i�1��HE��.Eɣ��J�F0È�XD���*~K����.�KI�p/�s�'��hWg���uw%S�Ǒ?�Щ����#
V4*8im� �ѓ�-Q�6-f4�˸q�T�/KC�=����$q���J�8f4�b8�T� ���V���N����ن�G��$�0D��'�r^��W��^(�VF�����:4|�W8����n��?�ڱf���~��*:��Ճ�N��{��+�8���V�H-	8��������xj��8`V�V�Rw�	�TC�Fq��B������9[�	j&��1��a3��IYf�ƕ
7��]5�e�T��?Q�y��7|�$��Tv<V��"�UB�L�;$��\�r(���`���8=��xx�]��WH\�ӄ9{��u���%��F�ET���kH�èFߞ�㍡w>�o���L�f]�r���EKp.����jFaq��J��
�!�#��������'B-eZ���.֤��c��*���)��� נ_�O�tv�>p���o�f?8b�9N.1��MUJӮ=>�n��#�)
?���ߖ���D�~�a�Ȁ��S�<�J�@�Ջ�k.S�gF7��2��LԷE��[p�������ff�;/{&Ip����!��"v����y�-x�B����h~�4�cO���� #>+�e�gO�ꎿ:��&�M�;nE]�D�xPfI.��pұ��0����#|�Mw���n�>3�N�ڄ�R�|).�H�o�������
��łs"9�[��Η�"u�Y�����~�Ł�
��P�^��e�������rlj�Hf5�y50�X�nV&~T�ǂ��6D���}hP�����"�yՀ����И���2������4WBL_Q��d��*�����{��� �b���[�oE��Kb���/(��j�4)"*c�}`�N#�ia*Sa��B�4>�!K:���u�6#����v���N�
P>+#E8z��1������Ћ�_��IG�[P���"�>�ҋJ�g��T�cAu�S�,u��F˕�!�҅=�֜%W���ɜY����������MxH0궾]Vg���V;ax>Q�	[���c`��nT3-��05��̈)'�g^�����z�/)����6�F�9�[c��X���)�]��4���\_�E�ܩ����Ub�X�k�Q��>m����a���jZ�����kWp\&f>��܏��¯9��̸�M�nuvy�\oaׂ����k6h4�2龜d�j�H��k�,qXY�@
Ƴ1�vļ����W�iR%S�MM/L�:!>y��I؎E�&u�)�T�J��s�ⶌK��F�AZQ�|�Ɂ���E�.fļ.�.?r{de5�י|>�ޤw�џH\*s�RW\���YS��F�7ʤ���ɛ!WbWTX��%�b���tu�.m�Oc������p�<��s��،#+D�>��-ȯ�
�,o����4�]�>�Q�:A���
�K�� �&�XA�x����;'L�,勱�p�!��/Խ�q����/5/g�X��X7�C{h�0ԕ?�I�b@���>fii����|�
���$�
Ll�Ç��� c����bs{�r&��[��`YҐ*�V���q��o��'�c[%�V����g��s�����ś�_��ə��%�\U�%hM�*������A{�xټoc�=��
Ib�)��ޱj��
3i�:#�S�6��i)&˓�r�8)ܬPN���C/�������@�����g�

i�
��J�o���\h��S���0B�j�o��@��%��4��t&i̩dJa����7�Mw�[� �kׅ�ڸ,ʩ�{�ۮ0��41�N�5{�m��ۀ0ۇ��C"���J��:�V˹�C=�4��b�]{'~	ou/(�E������H�3��Æ�+e|�t�
��PWîWf�)9�uT]���bh���k��aK�����v��ωZaʬYB���Z��9����8|�W�O�C<��UA*.�h��ō��7��t�ȇJ�u��>.�Ȅy���n�
oK��88�| ���!��K�G|��`i?g�������<Ǫ��-'"���\V9������f��a_�~^pt��tp[�)�+Y���W��$�9�4�"hV��<���u�W���d?���c���71e��Ep>�'~�y�j?�2t��D4vE�C�o�:4���K�޽����p��©������+��^�B����F�"�5�*c�E�UU`�O�0`���O�nI;;O����<8$CMc)N
]t'�Ė�פ2���Լo�?��S!n����GC�����hp���36M[X��h��M��'�#d�o���IB��M��j�3_e~�$}� ������[�x���=���}�q(sz��	�0���`�G�i4=s����޹c���@������Ԯ[�������꽼�9�)�������g0%J~I)E�dݱ��������#c��_7F�I��%��D85!�z|޴��v(�vg9��>�MЊϜZ�yx�5C�H(Q��a���m�|�	�i6�a�Wu��ڐ/�D���2���g�Z����y����z>HAK�,����Bm���'��Lˑ�\���Ӏ`��^BEPr���r�}�-A��"6j����:j����(Y6����?�o��(6Z�Fd�/�3�^DRZMT��|!>
�(�K?BP�6�u�����o��D�%q�G��+.P#`��uT$i���(�V����v�#��ܘ �"[��*�mJ��� 2�9��A�rp
��}����-�=�E}�&�i���}~�h�m�3�0��h<b�ks�����A?����`�B��"�ԝ!��}���z�@|TN�PH��9�əh�#��#ۼF}�3�v���_i���u�2���ܳOo���WEEE�ǹ����ۓ�V���RPH��P��CM3�%�^?7�oƸ� ���|�:��e��3�&��~w׷�M���/���W�LH$>�嚧�^�|?PZ�ML����O�c�;��4�IE�I�:�Ew�"٠*4u89�`j�������\(���5��%v>5ؤu}�Ghcj^�`N�9_F"ŕa6 E���[�k�N��*s�*��M�WjQ�?B�غ��A��WB����UAIl&T��:�W?c����
�l�;�R��OTO�R��,��1~���^'�{H�Z�&���מ��0oG���|a��3]�㉰�8t�i}�6���Ye��.��%�"��-.�� �0�t�K����,��:�<��^,V�Γ�My$�E�c��:	,��7rWµ�)����4J&�����������`��C䏏n_�;{��<��yb��0�����\�:&�p�SJN;@,�W8?�k�i�Q�c�{ �?�S�"�D_�>��K<4v�%��������f\�b�u�I�d�����.H�F(� k����?�O�T�_��<j);���;W,��vz���m�o����3a��ȷ6d>�~�ME��������$��PV�!�����zۍ5��3�s\Ur_v8$��Ex<���[�Ȃ\��}CZЧ.���Fg��2%X�To�&l0Wx����X ::�N�w�G�c�U�H/�6~�^�HU1|��������m��j��Wᠽ:���.0g���N����`�P��؁�a�׀�C���!b�J���	��p�I���z)1���<��Hc����
<{�ÄD�i	ܜp+`�;��;���?�@�7c����-��R��Ů	ݩ0z�?�9m|����_D-4}"�?�3�D��3f�k�Nh[V����c&���䅉y��v:!�b�K
�"u/U��Y���zE�t_���ܞ8K�ޚ�m7�����t&��3����&]Z�H����wA��%�
 �a6+�\D����\��h}�a�����B@F.[m�=�=X���0�I5���&_R��ң�@���&� ��8��;��+^���
!�XB\�|+���BM�OQ���Ͽ��u/�RAt�Ңa�SÆ?��d�wC�R�ޏ���]���>���������F7�����ƨ�̦�Y�ݲ����t_Жؚ�y@���㋐DI����U�m(;�;a������(�������`���={�R�
g�mg�E���縻�a�ƅ�FÄ�w�K�KϢǺ���kδ� �Z M���%����K�LP��������8xc1��vE�n6��b�����?�<9RW�|�m,CYj�2�$~�����a诪\�qx�Hʲޓ�<����i����M�X�災�7�ct�b;Q�hr�].59��2,��j����4
~�)�s^HN��?/�z��Y4,����_�jC�/���<*���!߉�~��v�ȋf�^��!,w���L� �U~U
���F�m��7؞�� r.+%��"�!�+�`�~�8�F��[��=u�T��t'	�#���~2{�n�Gkg�~����o,@��z�*pk�P��~��Dđ,G�X��Jb�w)��y�"=��L�b>a�,��/K�W��{T%���yQ�8����X���Y�Q�6�Sy-Q�Y�ڻKg�~[s6G��[��dQ��q�=>{�|`�����c�N��N�%�O�qt��P$��ǉ���xh��坹�8�`G����ޚ�M���T�Y�\q���y!�㎑d�\�R?\��Ó��~����a���L�A:���k¿�rK� mc~'!!��.9T�����.��D;ȏ/�O��b�NO+kc�oN��H���/�n,<C����6lSd��[�s89�2�c�'��Tb�dL�����s�~������+��"��"����+���v�3w����+�!�Q�ݨ�d�*߰P-~�͢�o��;��w����^kw�OI��j�B=�BP��iO).�f�)��� A�Hz:�i)�F۟��a|��֙�g��|xM� �_M��F*[�Oő1��Q���2A��~&;M3<W��wj'��V���`��(�~}��$Lͬx�`�0	h�n�2=w�����!n|���P`��ԄU3q��=��D�m�ʁ���(=3��kt��9T"�鮍/��t��N����ì=�f��J�)c�ɏ>
*���f��RV,�E��V�4Sz��&^1����4����֍\o�K�y8mU�i��FVb���0��[��.��h�Ǉ���~2M ?EGs&��ps#���Բ ��S X�`�KD�R=�?}���H���Hx�w�H�',��@�L�N����xB�X��_# !�	�[)N9�G�e��%�R�
�����N�cb��v�VU�>�/�u1U�ǓڟX�͜�7����IPc��B21�ɋp(�&gx�]T�H�������i)�ވ�p@ݩ52�R�n�LLȤE��HZ�9���B�,k{�ME�����r���xH3C���*LGKFդ(60��T�C�e�H���g���$_L{�3�m��1�2L�}��1�c��8�AD�F��b��AU�B&�^$^	/���
��z�;DUR���`d� E��x��f�>�S���z���.��a�0|�����!�<�������ˠ O^Y�@q�*���w�ce��Έ#� %���4�őBA�Z�e���g�IĎ�!lX*XAb���҃؃mDLDt��dU��}�$8>�E�#����l��-�Qh5Xy�����$��2��	}1�;��N���t�6+\����o)��^;F�˧c��H10�G��Bw`]8�A�_|�0��ۖw/ʒ	ߐ펄��:�?ϑD�����`�CTD^hs��z��2,1��J'�thH阺.A:F�L�32��N���ql~h�U���WF�M?#cl����Ge�nS���X_���7(�g�� �9�56��}�F���(Q�o��г�	t�]LJ	A4:�Fi�����4�ĳ<K���K!�ɥRH��R�{B���u;,�
Z"���'I��N4�c�ܮ��-�p-5]#�Ή�4�{�y,|:��I=��Q�A�T���ϞS��%����uU�z�B�qĂ�|��!��ް�A���(cx�4�i��%�jfE�&*m�h��$�h��_'�5�چ���g�v	L�3�n�A�~{L���97��, I$4��Y�£��~��ʊru�BI�yZS.<4���I[�\2�Oɨ6������}�j3��d��g�-���v����� "�m�����aY��o�z����3���c}R�J���=��tö%cFP�{]�Q!Nc�k��?>��=
�	�M�`�n@�Y�敶��L���;�=�J:΁�~�V�N�d�ݪd,cߊ�&�������?���q\�.	�8�n���Ӣ����j�W�w���?od�3�P��j0�xHP�H[����/�6"�R=@`͔%bN�����?i�U	�#w�ئ<��(<�[���"`C_	FimIF���iE���::�l���Q��	sKbb]�%VSр��=�;�ʬ�O�%U��&��/�v "���C�H��j��Eğ�-K�A��6�_-R���9h�߈��>���W�z�|�2|������(��}�G��u�y��8��?��V��f�È�;
��OEMknR��� PV�C*���N���v�|x����楉�_V�W��Q����s�0ef��N��}>Wo��(s�����Չi9� Ż�x6�웢�"������M�L�B��Q��W3�
�p>�_u{i�21Ɏ9��2��&mv �I��_i"���h������Tj��U���E�ș�O��}��fv���{�bd/�u������������d2f�~��������Vs�v�k[�}����,7� �y�yO�����D�K5��%�ba(N��Q��p��Z��_۶�Z�]����kX=��{9�Y�v����nQ�6t&Doq�X&v���Fj;��[{���E��j_Fz��(,?�M�["�5�ԋ��w����j;^x�?,�A��W/[�.�����r�������9
�ǅ�'Eu(������W��R�����
�xdݯ�ا�y�b���q��^i���v/vKZ���X�%f�"H��� ��[Z����Bj� �N]��o��p*5�7�Ͻ��P��뻳���(��U�{YS�0��؛���[��[h�O�9��T�֝dy��۠'�&z��5�^Rsb��5Rqi9n�+ޣ�j+n?6?���0�b�Vn/bB��|g�<��SG�Ë��ͷ���"F�t�;'�]��yt��l*�.�]�֮��Œu�ݩ� j��M�	�(d��ֈD��5��0U�Z�PDX4<'��A�p/L���H�J)�e}_J�	=�����TKDO>Q�.�ь��xп;ڶ,��n�J1�.�3�Trz�v±�B��F��L.��*}�w�����<��3b����e�/��!O�@-k�T��Z����-�����F���J�c��v �TB}+����r5j���c2rx�$vQ�!5^��v�w߮�xCM��vh:=;�+�=ا��=6�ժ�"2�HxmϮ��BO㐹+�+���N����O�?�	���G�*`��"�R����[��;�V�Vcg1�^
�����5�����|��.�Vxi4韥��}J���@���]�o�a|X�}���!�|?����̙���p7���`�3uuH�\`�,�>�ΜҶU�Abo�+�����Ӫ��s�J�I��r�����!W��WP�k��%��2�Yxmf�6��)�;9�^UUD�	�*�a�n�Qr#�{�����MN8K�w�ξ���l`��.�S���8��	��3\����r��2��ꔿ�� �3��hА`祚���Y���6���L�XV"3k)
N��.�V�
��J�z|�\���&���gY�q��aʫ�q�w���p��ŐǇ\C��n�fc�
v���⪦���pI��1FC�.��t�ޣD�d������s�/�c�ҼI}b��r��Ȩ�����k2�����U.[��Q���z +z�/�p�q��c���s����}���u�������l����f�٤��8��"��O{��o�a@f�6���	�����I�^�r��$?k�7��^2���"���ha�R��玧�I"�J��;;��o�����Ӈ�_w�������y�<\�_AIF �!��]C΂�!v:?:~�p��t��PE�Ƙ��o� ��æ�K}������q�Rn�5����ջ&=��
���D�xN�(���~��G�!�"�C�m/1�|~r^�6���Ɏ��tѺ��
��{ϣ=�;r�$̋��[�'��ِ�i�G�p�yN��#9�ҽ��;Q�!,�{l;P6���?S$�B�Έ7��J]qp��{�8Ch`&^���z���&T���ٳ����;�O��:L�8i��%#	�ׇH	$�a3i鲑Mꅓ�)k�t��s����u�- �#��FՌ��-
��.+!���|h�B�
��������9�DF�'QG3�����G��xDP₣�;��:�{Ѧ��纁C���S�6���� �xQ��u�^>+d-x)���e�G��]�{��X��� '��f����݂˫��h��uԼ��$�	O���YVL�ayt|�|��ѹ��Y���\�!���,�$t����]����ć�/1q{�c�������O�t�dj�vA�	�{�
�����8b'�O���#�
�o���*�B�;h�ET'<)K?(�-�_�?s�P��%|���-)���]����X��E���}u')��u"���Lu��g��OG����|�i�`1Q��	m���l�)ꖑ�������
�ӊD,:&�{�H���s2f�#'?kۊ�+g�*���~����Bd�)�%n���`:sI���32�����a?*������d�&�l����T�|q��ߛ05�����Ԙ@�q�gZS��M����?��7�U����9JR���	$Â����↬��Ï40�?�h��@��o���wg��zza�0�5��vN����/_P���Q���
 ��⒨�%��
Z�W[��(�
�;�џ}�2���EY�c�͍��d:S��"e�R<L�e�@[��DdgAf-H��3:�_���a�BCK�EZ��<Q4~�U>H��/>�3.�z&���/L��D�9���-��X��L��:kC��[�$�q���w&K_�s�6?�)���^bP���i��*�'�g�<��HL2}����UF���PIox�c/��\f���T	d�u�����\1�Ov��z`�da�FR�2|�'Z0�"�oR;fn���3�u7�2�A�+���b�kT�՗֐<�\����Y�$ơM������Y0��a�aL[���� Q�����j�5���ؘm|䃡�aX����{�슣VO�ڵR�?l!�1w��{�Z<q.x�,a,�EY�<����+��fP�����Aݝ�9Rh��Y����1�~	�.�^��Rs�'����0���D�q� |������q!.e�oY�_QѤ&�g*�J��������L����d1�>�(����|�up`C�`]�k]*���>��=��q]������޾����vz�Ƽ�H0��Nc�FQ�/���^��ܲ2mmw:J�?��\��!e���ϳ�q6��B�E�g��C�{��,�c�x䦗��2�8��@~Z�@<l�>�d�rg	.^#��<6���ġ\�7�s�0ww��L��|5��)�nq�kD�U@[,�	��9#���dКj��q��ȭF��eeq&��]HϘЁ��`���c(�H���ޡ��	�\��j�͟ɛ�5�F�ުR	¡H&(���@M���e�P�ș�I*Df���ޙ'��7�M�ί���o�給���g�~�Ukѐ�LBz/�kQ07v�:��1nē��U�nA��ymT�4��~�L�"����r�3���R�Q�����k��o��iˣk�H[T�����%���hR��ҭ��>�"���u~s�e� �JÜB� �[�_��/�&-�m�M=���P��4vL���2�+ķ��&7&
�@�e%:�XQ�����p�hD ٲH�����USȮAJR���q�84�S]}�AO�p+vQ�v3T�?�"�b�X�߫� eS��h1����������.G_˛�����uj�8�%h@5j�����(cu�K
��8a��`R+����I�<��D/Z��Q5�V�fC�k��鑏���X�{^���LO�ʁ6��o'f^5&W��;�X��IS�eIg�B&2l�̅�W�۔4��PP�l�u���i36;_cc���	�P���X��IK��F�ݺ4��5l��w%އ�o�tk�eM
$Cp�TC2�r��i�  K~�4���������iP�t{UP`�i��ٮ;�$a�J~�p�>[�(�D�[�i��~��n�j�Q�d��#�4̈́.$bWoo��>����� ���l�+��/�GُV���<a���.3�����s%�i!x�&Ey���]�;��Hy6�����We� �1��5u������ԃ� �p��U4�?(6�H��%]tV������Ϥ��9<���s��T�N�k>8C/A����Q�nl���2�O�10�-*A�	aH#�X�rHgΗj$�q���+�􋎤���K4Xx�f����{��O!�0:6&�w�)���� ��ry���h\*8@_4����o�����;���԰�����xJ�?����}�n+�𡂨x:i�>mP���Xp<-��/���[��"��,��!x]�>����?��pr��MI�d�t?|C�6T��;����s���1�h���D��q�]��	����"�mʉ��W\�3���@B�u�Au��Gme�k���.V��=��Hwj���7֖�!�U�\ͼG�TBrZj��})��p}h�jN���-����s��W!ݸ�$l��Fp����;�~r��A�l樄2j�O]��M��;��'�t�~����΁� -&�3a�.�x�[Z��(�*u��Pj��������-���o�WJ���fޘS˲��9AK[�u�6#��=�긇}1n0g���V!De:2�y�6ǂm=,b�*�d]�bJ�e�M��1�p�����/g@�(�X�<����'�Ϸ>�|_id�x��H,Q�O�! �:G*6'���xB�u=����_�k��,�f&Qw�B�u&-�F������b4�pI@?�����e�����f�YbGk�-�+�OG �O�����YO;~OJt�� ���C,��f�@0���Y<̤܇��;_4�@F��m�̒]{�#�����&F�x��>�;M���[�Q���o�ټ�~Pw��@,/>(���Ԏ$��o��Y(!�<4�l�vj(d���n\�zm���$2d+~��%"_#(��< Y�σ����J" �o�7����Ǣ~SL��Cd<�� ɱᶵ��t������՛U =>�|R�_8�ֻ�qv���K�%���� }W�n��v��0����e�b��eK0a��"rW�UkCQ��]���$D�W?�Ə��=���[�4do�3�G2.? ��G�9�ٓH�������v��7��O��^]�!�DG�K�9\���I��E���vuk�,�q�Q��D�
��޳��w�C�N�~��Ѫu���$E}S��������$(us1'o|��֯��=�����$">$u���.#W#�W��ާ�!W+���E�m��H������$��!l���#�f�#�6�t�MU����Nm@e��>]�1���H��͞.n�a��hX�$v,���[� vl�:�-�aY�H�������t��]QFR��*j!N-5��)�)�O�[Bm�Sŀ�c��l�%{�R_�<w�e^�B�<dٍ� �}#���It\�Ӏ�Se�?�a�,�U���R�m�����d��3�U��p�Ͱ�!E�밀�^���#ml\���'��IlX`���_R�`�6���E>9.nz3E|��K�z�\��+��V</�0�(9ik���z����b�f���l�lb��GP����lexQe��w����1���u�ba�]D�ny�M/U�WH4x˷'p�����OgG��ڕ���귃D��_7�Aϛ.�eu�]z��'sf��Uj:���T
�����g����R��Æ����E��^��t�<H��:����;�#W6#��nՓ���T����v~D&J���%A�2�J�R��B�߷��;�!_í�=/0�꣜�1��iP�z{��wշ\��\�>���պ&��!ƙB����}�焋�ӕZp+�rM2W�%���;�o�����>Ԕ����!�����<9��K���`��b�-��?R�-��Ӿ����aK����-/1`�t�u��b�ҙ�)���~�cq���e�}T�y��)�P��N�}�ĉ@Ղ�]Y���~��&�iw�O��r}g���ϘLX����"�K�6���vP�JT�N��C�uw)����x�f�5�!��d�����(�p񦒾p�-|�4�`n�Բ�mq�=�Rpc�ˎs�[�I���3Z�#�w �����5��/a���J����-�HM,7v��@�hߝ8�q8��nm�+<55'O�<��OgSG|!��\��e�~��پ�#������-T��EQ�_�3�p�q�����Z10.u�E�jKz�`��c?~�J!���gm��Mz��Z���V��"Jy��]|�}��e��8,_��3]ru8C�h�Ѻ���6w�P���#� Y���1q^��]�϶m�n�9�]�ɶ�ʶ�lۜj�亲k�w?Ͻ��|��^{�c�\���Q����>�Ǐ�[��SS,21��"�e.쒓����.��"�\�W
���a���J�>��������摘H�3x��zW�r�+���S��AS����^C5�2)6ג�U�#�O8�o��^m{��`L?�o�!�"�Yx^��=oG~��71��ح�6Y�;Z�p���>
}:�j8-�:��뫌��~��n=�F�4Ɵ.�]z��iBY>�W�w-x���P�p��O�.�K����^���!�Խ�Pӕ��P�M2���
���D
���7�"�Ps�3����≧�y���� �=0k�}��3!�ϖ%?��|�l��-����y}�A���g�)�y�M��n�>�I�t6��ly=y]����� ���:��^}~>7t����Wn��ӛ)�b!���^�]�ђb�E���D�5x��Ǚ�E#Y.����~Hm!���VTR6R�_����v7ҰE�o�&;�Ҳ��5�����胃ݽ�����f!^�H5�(�ư�a�E�L�t����Ѽ���=�w�#�p��Qy��]̷�hF#�vX��wڷu	ⵓ$���q�`��*0O%ۑ]V~)�uN'8���G����*I�~>'
���D�6���*a�o[<���]2����x�ҁ�	�ib����O���5M��|`|��p0�t���ܮE�� �L��s�����in��=��x�s` ~���(5�kH�uȖ��>E����i�e��k;ˬ�Ί��~�t����i-�� 5�g�����I)rZE3�"R���BU��\o�rIkK������0�Æ�D��;T�}��@)œ3��滏���Հ�3"���6o�T	�65�7D�mѕ�1N^�����r��7���	�6\�\i���<,'c.l��}zW�3�M ��|��Um%�B�T'hh	*|ǜ@���e���t���;�H�m�O��j���[=�b/���i5x����d�o�C���?0�p��c^>�Te�qگ��z߃-���绷x�5u*��`�S/WO��
�(��=e��T'Ių~�r��k	�?|�]I��`�T��t#�i��C�Hҿ�.���|�P��r�p[�i���\���I��X|c��<���*�%~T�/6o�hg�o��7j�6�:4��V�t��xTNQe��91l���no�!�DE���y���ž���"`G_Դ\�H~!`�º\�le��8��(���M��bu�����X��Z��m�׫����*��b)N��i o�ט8�;}�Z��Ta�ȅܑ�M�˚=^���k
o���&�jt~@F.60���psp���Z��)L�r�J*��QB��s��Uy��x���84��;#[�0���v[-��"�3��!r]��0�6p����.G����6�\��C5a�Jz��� ��_�]�u�Ϙ`�Bu3b�c���6|���������уj r�������U��0ȏ{Ͽb�OqYWC�R�aTW���Q�r��Eh�0UaI|'��I�kb^���,r�c�Ш�>��ؼ���l�(�cK��ăᅀV�b�^;�\�E@ȎV�d �:��OMr_�<#���^h�� ��F{/� �:��v�	���A�qõL�>b�3�@D�-���n09���:�n�)NS�ˀc"������ p�W}j"�5e3с (�Z�E	(�f���f?t/��˕B�FrM�'�@=�-��j	���ibVFSs��<��jy\�d����_�͓6b����,5	-JUo��i�@#^�x�D3t�ɮ��`����}4���V�AnV\K���3aM����O� /IŃQ5�9EF͢�9U8� ��`n]����� � $7-��U�A�K-;��F��ș��vF��e��g��tE��i+�͵��I�4�L��{�[g[�UU,5p3@vv$��Z��dR�� �"]"�y��71��^�U1��N�´/_aU� �(���xT�z�-6�Eh�G�"��䌉E~n�F�����nr�>,
�9e���#rT�؇�R CM��p�Q,z�8K6O�yn���މ����p�{$��v�=��[^��t��p�Im����J�,������̋�^E���.6v�3��-<Je��v�̋� �5�_�C���^�y<�hn�p��4�5 �_k^��h�/�	C��*�Y�Ԛ�u�����	����09c�2Gr�U���0�l�ւ0��<�L�E��fN ����W��19Q�X��3w&L6l���C
��̼K���lO��qFF�)OJ8�W%ov%Z3ݣ��0��	''�Y�@�wH���O��Pz,�힯�O�Z��/}<}O)S�H4%9ʎ>!*
���/��%�)�^N:D��&���n�+�?,�a�H�tEI�Hg8[�E�.Y	�I���S�}@>�e�����^l>��1��v�4�!���?�,�D��1�o֎:Iu�ª5��X��d�dZ��mt�.E���q�|�b��ҡIu��4�PV%[�FL%��~�B��dŰm3�g$Ӂ}n"w/=������]6�ف�w��}&�v66�ߎ�Qe(���9���GM:�s�G�W�BP��1��_�>�ZY����i�^)��zO/'0�J*�<��q/�<�U��z8����N&�7^���}��*�Ϧ�r�B�רR��M#����d5\j6�!/���?����"�)�c��F�@�7)�i�^�?8�ߛLdRV$�1��g�S�0�S��S�f�q�2�o@SxpLז}pLi�<4 �1��h����a��"�η�\�x;�v>qDU���/�\��8g�ζq/Hr �HaW�"��Q� ���,��t�Aǽ�F��?����˾��W�=5�QK���>2 b����G���J#�>�y�ZE�=���q� a+�/O�$]�ᐍ�#�шD8�XO�.��wzsJ-��X��h�R1m:�G�ުU3fO��À6v)<��v��P��Ϻ�Ԭ��)���̺��F����jN^(���]w�3������.��a��TX5���Ȗ{:v�A�V:D�,�_K�9�/͖K�w����kRY��E�lğ�iq�=�!2���jh�&�\�u�&�ˡTemt,k�H���^��A:��h}�<��f�I�Hx�T86�H9022h5y�:X���Q@S��B�<�$�V�1����H��6�V�K��"���}ME���'w�Icl�����u�Co���c}�հ;u}4U��9�	�KB1���#X�A���������yJ-۽�m_6�ת��@I� :�༤��u����s2���?����H�pHf����Eg_�L��-S)]|��&L�jFziІi@���H������]:�t2�_���C���U���������jJ�	�D���.��o���et7����QP�]�O������k{��Pc+]MP����7�%��^�2X�ga�t��52��hn�#&��#�O�uJhI�ɘ��0荚{��-<|S�͗��t4f��҉aѶ�|||ȺuY�o��Te����GC�,�k�t���G�0��ƈ[9��9�i���\�/j5m��`�k+�RA&���I������g��svg?D�~��U�圧���e7��/��KZ=�n�9�b����g��_v~�Hr�[��<�.}�4�oh�q��a#���/�f����D�=ԨŤ�%Zz���q�� �x��D��RR��H2��0u�=[�G��}�>�X|�V��n�o�x��q.�QQNI������(6=fw_��<g�B,~�~n����r���X�?y�p�Q��OW�׌��vZSnA��Oظ�E0˂�<W�H<N|BQ�'E���2����Ip����E/�n@���)N�����mϲ�|E�O���V �<��l+h�,�A��v6�.�3�������^�{^��e��r�������r�ъ���)���{�"�.T:�d������:^u>/�;��������!���@ȃ`I�.�M��̯!�`�3̜�D��~�X�����z[,
%#Y���@K+��M���*����Ȗ�ߍ��!��|������E�S�Ik�**�.6���'.�Iw����H����ߎVv��f>�����	��7#⇙8�6����e�4v��MV(Sڹ������1�rM����Ch�	���f� ��u?T���љ��q��P퀿�dn��:�+`<q��y���^��%�D'Js~�[�����C<|RL&��Y��g��#�i��	lS��QѮ�8�2�R��W՚�QRK�I
t.�$/��_�kD��2���������Gz�w"h,�Yd��Ml{�~�m������㻓&��a1&�2:]��Kg��\����|zx�B��=/����E�&`����L[4I7o�o"���Β��ӆd�z�TŮ�P`�����o�:?�x��\���� ���F�â�i��VSd#(���4���`(�Ĳ�n����E�H�_��d��h�}�s��V�=�	Mr�������Wc���>Z��Q��܊=���;�l<}`�8ͻy*_�ߝ�@m� fw��T�â4��Ua"��DS�ŘI?1н���^��1ư�K���H<B,�5�BˠB*W���ԉc��"��b�疌Ge֠�,��87�׫��O��2�u!�#x�@-v�E3�������PL�|�%6���!����Lu���u�����OC#$97�>`����n\�{������#y����F=P����/���fq�%&ʖ�7�*�i����	�`�mΡO��7)�`����ƚZ�A�(�K2ݥ��W[ㅅ �BNT�m$&7*��T�+���2tZ�|I!B�սƥNL7����I�t*U�Z)��3�F���*%���I*#�g"~�<�U�L�Li��B���e/������RgK�ݾ3kC�)x߶�#O��1�v�4M��C\�c��I�?�R�/�"BX'�X�fg(3_��a>'�d���X� �6�r	�D\w"��e�����\��dp�U�zȰ[�NM��C)*V/m�\LT�Q���ah[VF�������v/�F�{���Ys�X#xX���O��Į�|7>���~��������<�\��}� #(
E�C�#�یB�2�|�3اM0��[��4H`K)b�i���h�~����{1�|�l���]���t�:��/�~ΝO�n^��r�R`���n��HWVq����D��%����~OX���!"��5���,�v�]��#&��8aģ�>��J�c�dV��{��������E�C �;CWk��y�$�} ���q�� C�����	�@`5�ul-Ev�r����^�~~�0�E��:���X�|}F�2PM���T����Z��`yr,]�@p���Ⱦ@���E��z$-&�M���`��b�QZ'fc�Z��Oֺ��}����dI����CzRc{��=�"#k�'�y�C
�O�"as�*��;o$���ҹuq����E��YQ%F٣#�WCHU^e�c:}���k��Q�1,�v��1�$����F���'Ȟ�Y�uLуy�-�٧��[�G'Nk6A�^%��S����J���s��Q�[oD�U'j� N�^(�8��ls�Ǎ[�>Qy,��$O�$����c��:�s���a�@7�z�}Q�����7��`��$?(�X��l�jd�yzT�D<X��#vJ(�缄�m�mP����4����ДO�nጮ'@�^���<#�Qӛ��+���wA4���V���Q�8�V}� tu���[2�Lp�>�Db�bm�*i�m�x��'TW�6��w5GৌO�Y|��߼�$�U�Ej���W��T/-E��90�E��3I�$��/ZȼQ��߿��z@=�cʊJ��P�r@Tݐ)Fں���<c��|ɢLeZbI�Q����L5lH�h�@�b�W��Q���h���SH�$�V�ߵA�P�i{���xV&�@P�n0���:9���E�*�q9܂��o�&npS���٨��A�D]e�`n�\N �����jӊ�ػ������܊ޯގ����e#ȷ�W�'�nH\�oЁI	p~ ��.�82�\>c�蜜�{VBO.���k��C��9���v�|�y8QCI*E�%zS-B�s'V;�9�t c<J������i��Fz�?�w(�#���,u�@�L����?ZF��ғ@�fZ���m9���6���w֌�A	cx�B�)�6i��TcE���)��a)��M��1�w��
G�i,%D������f܆K�H?��,���� ����vf�<�<�l���M��XZt�R=9w�}5�hc������tF,��c��iVrrX��X,�Jt������	�12~�C��������O�����W�Zs$�5��)d����3��4�T�:�y!��CT��y�Ŭ10Ğ&��V���?�U[�4MEL���z���ԅ��Kpo:�"�%A�7{L�E'
{q_d�JE�40;u ������N�yˆ���'|JOe��-��,�)�j�./,{~�#�2��{����hp��~�&K{`z�k��"�#&▗/U
dD�e����"֖RG�FIA��K��
�5��Sf��Qg��k�����Q�*V�KfR��3�!h�H�h��;�Ue�|Ȥ.5�$+����z�שb�2S;/6ȑ����V�΢�V�Q C������Q"�,��v�l�K�z�jSZ�}�',�4��w��̤��s�Z~h��`�x��xUl@�1�Z�o���1	�+=���D�a&��G����9u�i�lS"�.\G��A���;O�q�\s�� �hSYk�&\F��x�\�ۅKU��Ͳ�0J�p6we�b�[��������@�q�(d6���+JWX4�������"�j��oT����%�1P[G���ٵX�~o��i��N��t��]����(&Cs/$�9�� �`�2H��k$^������[~�	Z7kR=_S���A�اD�&���U��/��Hq�R��6��\uD�N���K��� ��G��(r-�K !u��^Jp�S���8�^(9)b��9��g���V�Db�*�hvaڴ{
�@���?�4�!�#�cC��6�e���i3�!^�l?HL^��N���b�����������aQ�[�y�x�a�pָ�qM��-��VU�#4��a����TF�#������dԲGV�
��8�45Gն��ёΗ�\*�w]���?�S���EB�8��{�HSTz�Ďx���V'���f=.c�.zx�h���{��0�f�3��dYL-!��в��q���5xz�abeB�Q�/��ot�c�lJ]��K R;�`��l�"Q��Q�iR��^�F��ox��!���\��îh�*3Β�������N��;��w����=c��$��XKӱ&s�O}�rR�ij��I��*������;��:��(a|FᤥaمCռ�ϥ��%����C��!<Y�"��W 9�*�������6�j����e=��W	!s-�b��aӁ�3n/ݠ�?1spMs?+��iy;ᆭ�x���ѽJt���d�D��St7��"g(��u�P���u�D�3/
�װ;�9�Nl�S�V ���&$��Ju3F�٤�Hı:^,�/�!"�]ec���QN`7�6dSA�Xzkҥ���T_�l��+ZX⸺Ei�z4�tҼ��,b&��3��%M��Cr�j#�=o����Xk�� �X�O9ݓ44=Yqd��ܐy�f����!Sq![
��gt�~�H	�^sʋ�S2����%C�s�Xfz�	opq�+�e���9�|e�Hrͼz�SgJVK�MNSenk	�: ����p*I-s5��7�����T�,����ϰoG
�;SQ� �hS���}������m������.:��qo2�\�f��_r��p���hSE����%��M�8w�L��:L�l ̟q�玲`�3]b7G��葐��������gz��Jh�;g��	^Ű��hJsv�yx�l1��(y�@*� �^ [�g$����f<K�����0X	W�l��f��&.C��O��������U�p)G}\M;Xnu/}�z�KV�v��n�����X�ۃ$`;,����F �I�d�f�u���eN������t��4F�x�Tdtꊼ�a���E��y]p&J	�����Fӥ�I�ƙ���o���R-d�����d˲I?`�W��B"f�Z�UEuZJ��b`E�q`����Y�9�V0�f�8�:�e'K�;*�Ϡr�����;�2+Y�$�i���j;b[�6���-B����${m2�u W55��Ȓ31XSX�6�go�n|^A��mc�*M��1��u#B�!l���P)�P5{>&�jD��;�r�tOS����98�Q	�@(������K~�VV�>v^��Qv|���U����чj�1�c�����������@2�٪� �he�B�;*xU,oγ��8����.A9�<�5+�f|�n��x���3��Oo*w7!�?�T�o1�x26/�.a�Qe�"Xj�,�2����Ұ��7S����#1+U3�Q�
���������O���h0�Q�!��B*@"C+q��fH�\�ޠ�8"I��'����g7�2)s�܆���1$Z�*�р\�[�$��u$�m5����I��.�"7~��X[�n����82�N^�$d��n��� @��;����tǅ�5�{�2C�� c+��!����ϤV=w�v�^w�E]ש%�Oc�� �����8�O�����[��`�����/�|�t.�s�Y�$ld��o����Of��t�]���[��9#����h�(�&��ǯ��ID�q���ڞ������$ն�bP>�
N�M:��nJ�b�5�g-{�Ki��Ќ�Y`�K�$}����^oo�u���m`o({'���6�#�t_EfC>���^ˈ;�);�o�G�Jd�WF3f�DS�\ᨘ�b��݈�ϡ�w>��Gh�}�L�5����l~} �������S�4�[<N�V��b6���fY�J�o��h������`�oz����ܺ:ɕ)/��}Ƴf'�>��C<\�mkrF�_?y?��#P�\�Vm�@	l~��B1��C�������{3���#�Ă�����F�+&����K%��
1��ծ����a�]�'M/�4�F�Ū�{U�r��@[�W�#o��1�X]<y��״hRX
t�2�޷��P[�a������a+~.4�ٴN������b7i�d���4(A�Jpb��ɦ�GXm��c�u���Z�Tb�P�v���P���bV�e������w���pT��˖1X+(M�OPD` �X]7:�.����In���ם�q���n��޾g?�Z���YFG��o�z��]y��&��)jA5Ԯ\n�D�T9�{��gvJ�Uf�d��9pyx�p�۶�Y�i�oBY��_�lL|���!]��~zO��*�<C�>��M%3�_��A��=6��\�X���$ּ����E��̕?��w�,{^����4ojo��$�tu��}숌B��GQC	x^�C�~Ba�`^������ݾ:�Cm�z�j&�B��|��wF���u(����_�CT�7s���N�q��	���:L�*�|���+g(����n��.v�k���f��E�6_�ʄ�-�4���W������BQ}E&~��#1-R�W��0�����K^D�}yk�XUͲ�㘙n�H�g�ICo�B��^�q�}���Nڂ���~��Q����ɧA}�R�O��饩x[L���h��:��7v2n�S4^�������q&Q��[������8Uv��Q*%� :����B�6+Ol7���6n�|����7��d�����uc͞�y��d�%��V��<7�@��K�G1xHa\��轅�Z�����VOT�o�N��ӣ����C�7�� Q���=�SEֺaaE����[ܖ���up,�hB�d�o�x����ȩ���F���S����b��9��[뽄����(�r���T`���މ�l�d�ݎ��v�2_�a|�]��ͬ����\�r;��D;vb�t�	_C��)�HBԓ�%8>�:�d�<ɋ���GX�'VK��5m��r�YG`�����GR�C	�]�D��������ż��ܔt�������zN.����?��N�oE��%���1Jvo�	~�f���CBگ�i��j8�V��F���\����:h�r%{����D�,�!ӗ�{$h��m�!t6�S\#�l��I+�"�8���ꆅ}�a(1i&�������b�.�T˨��6�|q�Q��'M��o6s#�~K�sH��<4�6 ��3�Zm��'�{h((*(�~�]S�[��`�S�t'�����Tr�7Q�m�/{
�Tƕ8���;\��d��� б/�|���8�\�3^��ωϐn��/y�������)�/ɔFιҝŞ&�y�G�:�[Hkb���Q�����*���#@�!
#�x�;:a�L�J����	�˽1�AS;S��a�{,)���p�P�8����E$��Կ�N�(~b���YL��}**��'���@y�9�����>b���W��{�T�O�a�/o�|�����U�~_�^���t��B�[����Y�_�PM�_�ⵦ�L���W�e�s��5�.;�tX���d5�����E�i��\�|�v���0���(6�j_��m
V�n*/^����T�{�W�ɑi7�ӓ�+,G~%��D��dEAN���YB�s�,�B(��;�R<M���=]��M��I˽t�Rג�a�	�I�������~�?��;8���R=�K8��;�*)��i(x��G���%��mWpG"�?;�ƭs��m�!�� ��y[�=c��j�qߓ� (�|Q�j�PSz-!��_V�{��l��L�p#�_	mb�	]��ܛ��y���U��z+j,r��ҫ���9�Xx�TC>#V$��4v�E;�Y�����jG�M�H�,f�2K!P.[H�O����`�^�.��v��u��a�K��۔BN�
%N�k��UQmt b�N�r�Y��	�Wt��O\�Y�����X)@.fA�{..��rcǋ��2�h��{>~�#V�ۗ� �XL�5�)Q�pK���'�������BN^ŊR��}��~B�Z���cE�9�BT�e����I�^k�@āO���	|�;��S�o�3�^���ȅ�p����*?��>hзgba1-L�Y@cHC���)�D��қ/3o�נ)o�\1,���ک(���Z�pB�?�1hln ��z����x ���]����Nʩl�@8���`�Ȇ�R��,	?uV������\M��0���涄��3?��#�!�~p-��]̔Ɋ3�d!� ����[�N'���W��j߽���˜���uU�'g�z��7����Y7���;�u!��|�mIh���KF�G�U��°�\t��?���)c�&7o���5V2�)�#(1XD����qO���ۑ&
�x����ۯ�f�d�kP�~+m��1Sp�0�Nf����Ȫ_��zF_ZQ[��{���XW�%O�Ws�7c�0!ճJ�z����-�N "-��K-����Gfn^�v�I��P��O(��n�~�j��z�R����7��H����YsT��M���W�bϩ)�aU��� o �/�X!��,��3���zh_���%+�b��)'�By0$o�nz����?�Ӳۻ�I�$(�4��״�F��c�;+H�KvK�����C8���r7!��/��� a�MGy���Kp[b�J�J1���w4tm�j�x�'�}{!��л�h������?���ʵ���{c��$oKNy����㕚jF�Z��������֤o�%Λ5����#�E�@���:C��/MN�a���(��i���)�_��L�~l��Fu�Fl���3��L��/z$�]tƻ`�f�no�_e���YZ���N�[�5G�0�G_��T����n+U/BH��*Z�}M����=-��P�B),	�γ�k[��,��R��@�-�K�m�9A��廫��g�)�"/�OM�)��]D�h/`D�3�K¡퓖I��-�¤��Zr_,�7�\�^����FL�����]`Rݶ�"�0�����������#�������gQ�~����Z�����-իN��>�'���ş��4�?�Z�8CK�qh��8���2�������	VFfd��^��#(د���n�S[�֠<�)��%��ʯ ��7k.��n�uV�*D�f�4���t���`ٕ�P�*�8�',��Y>��%�i�5��i0l���.����)i8+i,��%~�+^����+b�3�E.����&϶��!�@<�>oC���0sjQ�W�_���#4�NgqP7<R���2�X�(.+Ã ��Q�]w��{�=.F�f�9�0O�d�)���V��VP��y^�*����;D����b�&�U�˥RC���{���L�v}�#�؉�#������>��5�(!ձ�h|kBZ+�B���Ò��6�-�/�����KU2�Fa� �ʲ��JH�r���j`4��U8a:ucm�|�Q�V�U�;~a��<X��d�z�ǊI�S����v�����$�6,0�g�^IF���U�m�Vcd�/s%?�!��ǣK��3�H�hj��&�������^�K�n��P��#��c=O��_�L?=�yY!�5�\R�߳K�:��3H^�/0e�������������)e��+��&��F��Kh5�k����5���9���*n�^�r3��J��"�݌�����2�h����c��j@4�Id�ʶ��ݘ_g�� ��L]��)	�E7�L�r�xb6rX:��YΑ���}�Z	y,K��-Ag�^Ɛ��j%��4m��j�V�SSR@�p�/=��zʔ���cT�	}\a.h.N�����;�C����6HH9Ip�s����,Ӛ��ٙ`��P��J��8����}�o�����I�Jէ���a��Z$�ױ�W尪R�>J�*L@=��
;����z�6l�GO�o�j�d�F���mќTK�j2�Qa�����C���q8�j�QD�6���t�%m� �E������.s)A~a	�,��|;�Lu[�`_�Nt�-n����M�ߦ����>K@<*Jn�D����5�z��^��I���f�4VJ��A8.�(Z6��h�.m]���.��+%�2E�2[� ��+@&�M'KW���ת�v�[�|&%Pp�Qꭟ Y���#U��'�m�,'�K�9�"s�h�ι��mB��2�.��9�����V���u��:�F�{�#��O1�B�����}��&��<�j0��QB��i�2|�D��RV�9 !}U�A$[�&#�MN<���-�\�bS��E����Xʊn�w�Ag��C�|ki�zD�2\���9|K��D��T�h&!���D�:�-���Ss�IC�����eE�{i���Xg��,!�ա��Mlԥ|劬!O��>�\�}�|�e��e�\��Y6W.�B��-�͛��a�i���u�����M��m�P+�{�nSCm7�|q����g�6���H��n�Ek����K�Pj��:�Jܜ^�J9��d3��\WQ���1���ӆ�GGq�Y�gPU���R���p�J}���t�o1���"�Ϡ��GS��(l+��+���7�ZD��J�Ax�s.&�'=n��W�]�=��Jxa,�I�]-	.��!H���T�E �8�8tMl�������FZP��%�OI-�Ѿ��6��<���6�����ߙ�M�cz��1�wn(
Y���ԟ?kQ�2d=�m|�"^�zʪ��=~�%����!{�L�]n�a�U�ʥ��i����&�.�p�u�P��pH�\��(��I<5Ď�ns'���e��q���õPbP�T�n��fi����J4~����\���!�=��?�$욉��n2- �s�Yj ��`����0w�F�ֿ�&��dIO��ʆ*M2PTa�f�S`�K�;���&IB�ۅ�*�+��Wb��K��٫�`̔.�U,p��"԰s
�i�J:7���&�򘎛m���i���u検��6��2���o�;��*+��E�8SR�Ԧ-�Z��cųS�dG%�]��`�U���C�Dt���^�������>���$��~��|^��s�F�o=(۽����!�&�.*���"�R�h����;=�a����m�a(�@��q�TU؏=�z���F[o�&��o!�3��pl�Bt�����4��aywխкȔb��
�"�p��x�T ;ϙ����"�/&h�%O�Ϸ1'���<���<�A]�F�)��Kl� d"!.fZh]K��8vH��.�-og�n���UO[d��z��Q�Vq�֝�C*NUS��nRH�M��h�7� bu�,�E&W�^� o*���;�(��ZI]Pİ��|7|B�x���N��B�kVJ1o��G���b��wgT���wi���y��IW�B#v����5 Z�1F�Qͻ�;q� /I��#R�)҄j��ʗ�;�q�v_5�Ӿ	��8~�!P/������F��K�H�?uc�$��H��؟��5�m�F�Wܱ(��F�2�h&�H�{��Υ�jG�r '],���T?�e~bLe���YH��%����N�1o��mq�	����A+<�!.+r�a.:�ui�E
G,�������(����,O�S��P
�����<B�a���j*��O44s�n�pM8Կ&_
\��f�p%�2%����s^Q���:a4Z-�wLT�\�3������|_�Q�h�k��#K6F=�����u�|��{	��}Q�^z�G+
�8��a��m���VP�w(,dD����� �?�O2���5+��q	��∖��&�:�rRj�!�*��� B�O����|qd��Bp����SFt	Y��mgD>�H?�zޞTB�� 4#N�p�j�Փ���m��'wȷ�-����q�8�g��ׅ��^���<�0:0����G� �z�$>P�8��JS��o���^X��	0������w�> �U�j<Ɇ$�ݍEW�hj�����L5��Ǐ�bU�C�l�r�yο&#덢."0�����!jV�)m�.7��Y�B���[eu˩��!�
J�rX��w��������/8��(a����Aa��7�PG��	������pdr�G�'��6�5�����$a���1���$P�`�.gp?�Y̯?��,ĉI�(@���?6��)���=���^�H²�6*�VP�;��	?6���B$���n�w:Ntz������d���$�ip��]�ު���z��w�)��X�IA�m�0�ri-0�*�;���]��7��(��%)�0J��b1H��G2t��D�)x{7K��#}VQ�K���G���pL��MRii�I3�4��\]���N��v�я�A#��%����ƿ�u����߿+�'�հ%�&|�)�
%�bV�C�t1:�(m�ϟ�Yێ�;�ZU��D�v��5�ۅ�؈�"7tc�:';�r}oW2�
$:��	�,	L�E>3Ǖڷ^����\��O�C{�O�`�q<0�2�9�&^`J�仲t�(� ��:��oH[DH>�m��^�����jd�����z�˴H3|�vMɊu$���V��
Cm��AA�r�@_�'t�<�vv�"� �N]F~����GNP�����ˋ
 ����H��{�U���)��U'!o�O�����a�|�_@z�U~�R?%�Z>�xn�缉:�*���j��p��>�:�= ��Hw�$2�k�@�U��hQS`3��?x��ڿ�N�������p�Ǩr��f�������mߛ�|a�˅0��{$�\�@�_����wU�`�Z�rw���e�o/�	#�m�����3G���wޯ%����\�������TD�?��o���Y:�>���[W<��Ewfu����B�~�<���Q�:3�	�؍���<�sz�z�nX�0E�{	����(��l'b�pxu&���)epw����Sϕ@ޣ���yn�les��Az���*�V�*�No�wh�(��f��N�2����k�N�˷G�������e@����6�:��k7Ɋm۶mkŶm'+�m4l�4���h�h�6~���]���z��Ϝ$�ȁ퓎)4�EX�Θya�rc� �4�>�d���be
�_޻+)�'��q8���Pӗ-�Q��D���ŧkn%1Ӭ�0�_���8�֎]!^�#�ވ�-���YG*���l�3��o�X��Xh���Le�]�;��pN4G�M��-ۈ���+G8
��&%�	�j�W��l�C�_N�`���$�bn�3H����>��l:���o��b��"����,}X�aXԡ��(��"��2�6VeS2{g�-�+D�Ȫ��|�n�/%+ϫ܂Ą��B!�dq���b��Q�������_��(�%�胥�;}���H%e���
LR�Εp?������uK;�z��A��y
h��:N|�s�B�y�� �=s��~\���~� ��90v�6�:Sʊ�СR`�������W�V�n3Lc*�.�K�_m�Iv�������Q{�]�E\�ڌ���y�I������QE	���JU(=L�Ke=���g�{�G�{�7��d��� �0���yB͉0�/�dJ�+k�C���;����J�����7+�`3ZzW���J��k�Q%�h�t�;.��VT΀'�1��W��p��@�����s|~�|�?=��]�ӌ����4�;����"a�4�)7�ǅs��N���������ݕeDç\�,�^gJj`A{|��(�>���w�ǩ��"*�pF;�l�Y����n6�!χ��R�/2�� �p,�X��_�����]C(Ҿ�V��#��dW��__9�ɒ-I�ţ��q�K.�v'�E 2ڎ���u�@�T~%��5N�����k�dy�m}t������nH{�G���Ƕ�Mn����A>��	u�~��%����f�gK���
F����r���gՙ�f�}ø�,U�$����p(��#V�	�)#�9�ФNKW���GlZPu���qv�ו�^'��nPO5E�ۜ��u6�T�F�R�:�� ��(��qB��f�Q+�Z�j�;���{&Q�}�hQ�A^Z'�jk4 ,�1|���*�c� �1s
�dR�_�rv�������4��$�n���ir�!�=.�a��$A˓$A��<���w�w��=3	(��C�^�Hf�J�E�k�����L�,�4�Q��f^���Z�%PTs\fe����D���x�'�����o��<|�����v�wЉrsC�?a����ώ�4��⪼GP"����43���a��)Tb8%I�/m�,�M.�ܖ�rdt�܂��a�5�OZcN(��~�k���n�Z��A�e��e�̭��^0ci�c���u���H&@��9�m�:��Bq���ߘ"�2��K��	����ϑ!�@oUF�Na��̕2�����*#��ˢ#�6[O�` 3t�w��������$xV�� ��%�RE�{��$���)Z� q��M%�����d��/�{����c�>��Ha)*��o����|ʞG;B�Q���βtB�sH�%N�v� ��:����h����Rip�ө�m�H���,Uf�3 ;	Կٶ�R��A�W%�*�$[!Va��.�>���γ��B�@�	j��*L$e�jc~2WA#�R����H� ��z�(�����d�Us���o�g%b�E33i��,&]B�\������Ԫ��h�gr4�e��#�aưT��	�ҳ�;�m�Cg.d��ر����S�~���O�_�{8+�LvƌK�sz��¸8�+^�u���ӭ�'t�hC=��(�X���{u/w@��kf�ʄ=m��IF��y�x���Q���&D�
gP�C�4;h�*���^$�Y���/�1{K#�\*:��c)5�u%�IU{�_X�N<_{r�����1r#��������uƛbc��0Y�x��\��9��"7|�g��:ʨ2M7��Z˘M~�v5\$B�M�y��5��3;��s�(wێf�Q�Ԋց����e>c�|\���jR��.5�`�C䳒aC���'�'�{c��O�w5�.��B2l
�F,f%����wy�=[b�jX�͝B�g�ܘ"٣s�2Ft�[O�A*_�O1�U�i��Hp�a�'�&�ѧ��*��o�ۅهoMP��l�l3��`����7$.h��Q*^�;�i*���_w,���d
}4Hy�9c��db�&efB��Ӵx��z�5� ^ڶ.�� �D~�_*1���/�%Ƕh)A�^l�����̢T�O�}�+��O5�}�t򔻀-E�p��O���_�3�9�
*$t���eXB��S��S#p���tF1@�Pytʆ�:t5�=/J���sٱ�[G3�f[e���������J��2�@���H�b��/�W���F)w͇)���/5�6�s��'_в�'��~S��㊵��8J�#�ژ��98Dl���F��sZ�ۣ �V�ŀ]�������:jh<��K�D�ʺ� �EA���Β[넚�9h���
� 8Zg=6�?h��C~;���f5����3K^����!�+�c=�9rxN-ޠz��x)Er��~�+t(o�:�E%�oE���@&5^�!��������������/o�4�_��k����� ^dG"��Tb՚SP,�q@.��f�2|v"�n�À�C�v��R��̀M�-�l��󲄱�hݼ��	l5ٟa��`����g�S�3�
#?�9����@��8�G�&�mѥ��,͌w�Rl�bl!��!Uj�(��t��G�G�'�d��ĝ� γYH8M��N�%)����]�b�ᵈ�Ϙ��qwI�(J�@Z�^�����|w�����m$���t~?��E�R���8��;����úM��n\å��7`jX�eO8C��� ~;;R|6	�,~����Ǡ+P@|��xM`}�X_M���9<�[�c������Sd����M �ݠy��^>)Epa��y6�,��6�Np.�t�a�M�
�a�3���,Qz�RM��`gױD\m?��XS��Qn0}�g�J>?G0.S��h�<�L�9�`�D��	s���0ϣ.��E5��x櫶]��T3��/�	(2Z
�:I��x.�f�l_i�}�F���L�Q�����Z���|s�^��!�ߞ�8�L��SF'�����Ʒ�=��v�:�������n�&�x�:�(�P����������|AgV��a񶢸�E����|��|wi�����~mŁ�g�8M�ā�{!,bu:8j�	b�Z��scȹu����i��z4�e4&5O�_���D�	��]��̈Lˬ�����wL+���(!�ݰ��οj�c�[Z�鑌���T���W��7J��FWn��j��ov��R��Vؓ�Seh��>�W�۴��'	�ژ!���g����ЮP��ڛېO�*#�˗���1\���[�%H���ˋ�f��Ȭ��=�������E	�s4���%�\'�Ϩ}�Q.�=:� 
��\Ku*��r�$��M|-�����/Y��+���
���{��P���N����'΃�K�X,*G������E��ۨ��)��t����z��e�NB`�硎쫚,v�C뺊��M��XMH�m�L�pdh�N�Б���'G�ʅ *%�	�#�W믔��	�w��곫6�f�X�����k���%��f�m�*�r~E�sWV���s�1�H{����z����͘<���l���ŔׇjFu��i�fL�`�\"�˸���O�G"��Ɇ.��������R��U�� �������@�=�#�]��#�wG��1H���^�˧�G�����u�"O��$XU$dHc��Х�����I�-�N}���X=���Tqpwofvv��%6{�����I0��쐆`1�����t����^�W咍��Z0�~�[�e�`��8'>R���%K�!�׭o��R��}��зY��]�<}������*B�<]!�g�_I2�KU�K�gKwl���b�-�W:O������{����d��H��}���o�4+{��^��b������Ju����|�׾N�u�Q�3�5\?���,JA��b�%�!7R�	Rn�~JDc��}	����ia$��Ӳ�:����[ai�"Py��I��i���`Qʔ�e5c�@�n���w�Z�l�1�P��ch���;��= 3��T��:s�3���W���7�H�m͑(��Q��U�Hȶ�hQ����s}��x&�`�+g�W�8'���W���2p�Ce��� c�LQ��O~x��R��ےGޒ�5����ʭ�����H�8���]�0�_U������;ib�&�U�	�3N��'3p�]Y��4#��'�]�7X��-�^Z׿�/U8�.Kt��$y�������K]v2I�]R6Z���� ����C4z��o9���{�u4J��X/�v9ú�y��g @o�z��dA}�8M:�g�� qu  7��-d�J$HPۅ������(6�UXz�����}ރ�350J��Ν�#�5~�^��o(i��u�k��
��?5��Ώ�Ck�rک�y-xX�4	R9��	8�x�֙u���H��lZIRe�G��)�}1��W���v���Y����MΔ"?U�U������C �k�pY4��*)�9��6�'�Ͻ�8E~����ҿ��4T�Ӗ��zc�%4��!"~
6�;�h[�<!�u���0#��.�G��-�z&Y��r-��~���ܶ�Y=�����jp���I {h�fe��U��8_�s�X�a�}2�f�&~Uq�Q�zh���~�r�eA���/T3��P 2�m�G|]�ꍯh��Ɛ|>; ��6+�i�-�q��Ġ
�B��S"�}j���3<g�w����!�G�q&�D�Ue��dqh��32�l[�2��~��B�b� ౨fA�.��Ӧhȴ?�U4ҝ�$e�x���d�n0�6�Lk)��ˁs��/�kK6a���B���^W���w�R���Y��yq�}�WM�y:V2���ZF7`Au����^u��EgR�rQ.k���_���*�wV�["P�ҿ'�J��5�W�&��~�e�M�������O�v��B҈�vd�Y'��t�ո���!���@ԙ�'�����n��s��7�s>��'�����T
�B���Tx��dRqz��	oD�� ;o�Q�a5d^˱�d�Z(q��_󆻩��S�xH�
�y����Ņ�#,����U�Y���:�!�y��*���u�Ag�W�G�W��x��J��|\�W*�)�.Ϡ�� b�a��1�"���nw#����,��jìۄ}�r�(��Y�x�o���jm�<ŏi�l[�Oޞ}�o���N�W�V�4ƌE�SG-�l�v�����4�<)��>�@��h��[�����*�eX��*Xw�
f���!�W
Զ�ԙ+�^�>ܨ{��P��u"th�?��	;G���ic�i"Y86Q�@�kl��Vy�[���%q�
*xJ9�CN�n���'��+Ͳ皂b�wc�/�I�5���i�{�{�)���\�jc\MhEK��VT6w�mSF�c���I�G���U�1�c�vT�<�1`}-�rf�b�4��Zܖ���O�$,�lW���L6l`%B��� �.}�kA�c7ɜL׾*4j�X]�j��B_����x*�h���S]�����~$cQ0�� .�o���l�z8]�.�+P5�.IU���]��a5��&�2��ৼ%�q��-�0���̉��
zR��l,z��5U�e�RP6�˼~����5J�܅_"��=I/� �#�P��6Ϫ�K[�7��e�)P���2u' �X��_�G�f�I�aSعlh����!bm����LW�b�g͍p�ù�'��Q�kt��oF9+N�$�(�A�0���;qr�B�y[�Ԓ��.�Y'������Z�*<Js>d�y���d	��`[��'�P���(��wBM�>w��M��[�6<!9��V��ѕ���q0ɏ��'o�2���Z�l�U6��������j�*��P��q�͖��z3-pX|j�=�օ���;,������^�-��)�-&r U ji��$]�^�%$�Z�{���A0�~��Z�B>��\�/u��3���^��MQ��д�;ܘ?U�ȼ f�J�^
u��Rr�{�s&E:j�9�\�;���G�P�ui����X
�	3���8"�����+�|J��G	he�f�/��z,�UX@ �K@bڽ�`��,6�j!�>�mP�w��I�׼~���A��}�$�T�h���_��d%��S�a����� �Qϳ�]F[�/s}�)~Y�1��c���T#��Ā�P��*���h����,�J�z�غ�4�;p^D�<��ʾ�Ok���H��?(�[6lC�d	�y�$э���ѱ|�(�
ŦRs�y&�9���g)��m�*��l\L�]bο��H����]�V$����vt/���G�w� ��\��{�WY��O%���!��ɵ�sU�,Z��%gY�@�0�577�1 ���Xq
9���2O�-��m<4��� �4ŕ�����1֗�}D��P�G�ry�f;sZ-0��ƴ����ܗ�w�8�+%�.	`�Bw�˽fE�~�u����a[0J
}����ta}��m%�C�8� TG4����a�7�SD�(���$��e���eSc�r�VJ�7�Jo����ë� "B�"�'�"2���Ӳ�"�%∃�j��7���M�e4����e�7l��m��G�-5��ݰ���tk	��G�E�A;6V�yI�*}4������t�g��M�VOi�}���Bu�'Ն�q��'�]���H 7���Ӓ��hd��煝#g���y�T>{��&���e�ʁ�J1�{i̓�,v�b�6n>GO�����ⰱ_>����S��g��դ�Z;]ۉ�S#�}�~����O���G�˅	� �:�(LQ���+jU���>�-k3}׮%/�M7G��4��7�d���D�D�aת����(L�S���Hѻi���^X�҇�I$��]J�5J��f%�m�JO]�e�U�� �d���n�̱N�s��֝;R����M/�F�hP����L�i2�{���6_�S�Y1cP5�_��P�[�eZkTlxt��V"�_�:������1e14���IVO+��?��x�i���P�}��B���p+�{�璿i-$w�5~2�؇$���K
��:K��.E
���xdBt¸�K�)�ߺ#ޙ�ɚ�����e.�%��^�~���mǵ��G�m�S�آ���6���'��C�Z���	���e�EP��2,�x�}|ۊ�p�C��'�[鷐��K���K"�b~/���b=ʯRl421�P*L�*���	�u�ɫ���ޙ��L(D<S�m����ڑ�˾��n��S� ��ƀ�{��	�f��U��K�O�K_��X��(�2[\�v�]4��MN8���;�/������(iiϒ<iL�'$���MU:��J g.W����{5��7�}y�_f�˾]�Ӻ"&�>���r�O2��~%�jH¤���s���3Y�:����9!\4��7��S�{��)�f�]r���4c�s ØD��n�d��H%F���j�t
ذ���&�Qx=�*���~M�l�h�V�3~	�y�M�a�p26�i�虞D!l���O�8�᱔���0���]m��1�ER�BMy�����dǝen�$���N����86�¤�hؾ����2�8��|LA�h�C�%�M�3H�L%�m�6r��[��e�Pwӛ�Ӌ����Y]�o�K�hs�37�����M��)Ц�2)��슋�+�n���|�m�c�u��;���)@��"dbK�T|�~`��+<m�����,��A���j�Fk�{�(��z��U*�;�1��"u����H�}
1G��͠������͂We�����ڱ_�9;��@�dk��z��;��uak��Y��ŕ���:�f�|!g&��[@�M���S�S�~$6k�2��ƌ�����m�>�a#��TR�[�8j7�.`�RI�gAo��[��޸�����.,хqY�~��bΉ̛-A�e4U*��_���R,Y�9�+=Gs0����'�+"N���¨�~J��9�X�,Eyz�S(ڨ��zb)m��ʸ���]�ojf&.�9s����I�0P�d4��۰Ş�}�E��U�����7c�􊳿�_��6u ��حW��Ȋ$�*~~xSt�����g�NN*̗�7^��K;�;�9KY)F�"���#��X��*;A�����B,�+��z��[!�`A���kp6~:(�;��c��(Ǹ�iè�k�����k�l���V�Y$���{�<�|u����=E_�GI1e�kT�A+ͱ]A7�7�1����`�F�/�c�3�ryd��V?�P�˞��˴��l���������';t��7��5����9�p��6��hȲu8~����$3��2�#��t��w�6�1��.�y��oʤW���Α�0Z))���]B~�C����TL��M�*�lvv�6�ڏ��z!1&f%�Լr&�&��lGξ��^O����jA����0�VBx��آ-�rX��]�((wt�3L�H��I�Q��~Յ��^�w�x`�n\�{��W� �&Q��4�F��<�[�y���F���!��
�5�3�
��Kq���R�An�إ*���X�{�"�9*�<��eA��e\�i�l��룛c�`��Q@�r؊��˵RG�sp�ø�&i0
�)��y��^�I"b�3��h:��4�\z�V�����!v&�j�Q��ԑ)A��+�t؇������|����\�R}�`�񟶤}�g���a���F�k��$�9	�,�Cv��C�t��V���L�nN�̘S����M�%� ���yxS��D���_F��}�퉴�哾�c�c����-�j@����f4RX��H��9�)wl9�=$"�E���}^`��MW��[,�R�_��"H�PV��@��JR��^�!��4�k�g����a��F�q�i'��78Ǣ��c���ስ�|�eZ���#^��8�^ 5�((J�!ٓ%ޓG�^q�SP̐r̸y��A�=�r�7����{`���D�K��3[�����T�W0�K)��p��y����'����	h����΋�#�3P��EL�K�R���8��6Q����@��Ӄ���ӫ�ߥS;5�K=n�r�G���9�5�P-}�zpk�V�S���O��yg0-�D�!x}�{����S,�ģ�������jx~:��>����q6��d�F��Ń�Q���]��x�h�U�~[�-��>�5��2؎
ݢ~�4�i�f�kx&x���s��\)}%4�>j��Af�W�zT�!�4��,O����!�q�a��e`�3aVh�	���HO���kbi'��K5�vX6%�4�Ă�bʗ��+g�]�8S��Y�v��$z�E�:�~��m��`?08�,*�x�]6[�ȩ��N�H�9O�J:�s�c�*ǌ�!�RːxRSy�G������'
�C�@�A��@��G�j�!
3=Wg�o��@{M���R�s��7�d+��6�&8A\��?4rѤ��$]�����$=�-5K�ɋ9s��xo`�w�}v4U���'������Vg_���*.�;�Px�ѭT�j��L��csU����X19}���C�$�ome��t�ǋ��j�N�������T没w��7Rߥ�a���w��3�i2�N�͙�N~�|Z���X!;��C���r���)J���Ym�Br��
�rOD���3 Y��!���5����L�����2�z�AP��FT���F��T8P�,��Z��w�M��:
D'�ڝk��h+�$Q�g:�+D��CK�ER-�0du)l�1:+���WEAZ{|~֐��ªO�)@�&�-������蓕�=,d�2%*�
j(��s3<$��������w��ʸ.}xѷt�0��f�h��hQ�jY��QL>_[R����3��w��b3Q�:�xzc,f�*�b���Oន#wo�ڀ[��4�t�Y[v$צ�6�� ���(r�2�����(��^I��[�چ^�[Y�_��ﲺQ� �H���r�]BH��%������bv�%إFd6xs�>ͳ����0ߦ��MxF�:,cQ�>�ے� �x��9q���So�;�=w���|j�%�����Z�7bA�d�W�H&bNl�&��S.�x�Lyا| �G�l�W�3c�����Q�eB�
ݚn�_�n����@A@y��h�ԗ,V�����_��|�@���8�s���h�^%����<���Y��U*���{9q����0+KCUQ�(��c�;��!�I����/B������t�z�8�u�$�ON�z�j)��4ѐ%����)%�zB�j;!b�ݖk�/�{^9z}s��%~x�t}�
{k&â�i!0D{��,UĕK!_0V�o��:��?�f;�o�.*�nY[`�ĩ����0	�W߲`{_�����}��/{!|�H�_\Ȥg���t���D����ɼ.ڙc4`��>�q�t�ܸ��w�Iƛ����>ȱ�Mj���K�?'츛��c��b��%s��N�`^^Jy��f�c-�:�$o�cg*`s"��zm���Z$��*���Y����j��wAǓ��W�=�L?�&q��.��D��Ȱ���a��]���1�x��k�J���FEɹ��-R�b����S)�Ck�5fvZ�c�Me���4���v�{��k����a!���,eU*��-�G"��r�TM��5X�~,w��p���@|eG��[X[��X��e�5��u+�|�i����ܗ��c��:�Pv����D���]�����Y*�[�Nve�C�q�[�c�h�"���9�m]�]�#bl�G�VL�����]��	�R1�66��8I�(����(6�-N��Ro���������r�`ށ	����Bl	�b�I�E_M�^^��ԏ��٠V�� +����#�5D��_U��D�G�����i.�i��S26�7Sg��nJ^���Ba*g6-5_�Dbz�
t�'	���h���D�L�����q�����0�/�}g{N�OZ����T0/na��K����;��㧷��M�)O�@�蕯�}o.�0��B�g��:J��&�+�FE6<��%0T?�6�DG�(��@\i�VY��/<��*of�S<I�=�.�<&�z�L�g.[���+d�'��>%���Q�>�&�'�����"�}Ǯ�y��h���9��*���1AB���.�!�[_r�y94��AWo�����������)_�Ϛ�6O��rB�p���i�o��d;��X	,,l�n�.P��i��1�5��j%L6H��uX�@MɈ
��@�W|l����E��cs�4��:5c�)pU��`n��x�p�G0�ZTۤL��ж*-�����9T�b,~� x���\������~���7�M�Ȧ���DP(g����
�bQ�~��,d��Q�Z�z���(1Ba�NM�v>��%"Cl�2,���iX&&��X��D&�v&�l��<q8-��v�+_����y�gB�J��D$ )��-�t8E!� �VA m�Vb�d:�D�O s5���A '��T$������\8FSX�%d?�H��F<�1��� \ܛ�vA�n"f���~)�Z�v������3��d��@���UÂY^�����Ґ�sT�
�\�ղ�*�(9��bk<�-hٮwkrk�^�{y�����lz�h
�'��U���W�&����?��/p�ʴnM��+7����oMpI�oU9����3CH5x�M�L�,�\�ј��K!�s��I��j��|���_	`�=I���HB�Lu�M�{\��UHc��fד������'`��(�y�F˨�g6�D�����Y��|�d_ϕmhD}��PPD�i�h�%`��FM7_�^����V	��t�;V8�aĴHFii �4IU()�����B:Ү�IoL��QK��<R����T�%2	�
�Whe~Ŀ���f `{6Cvf�RK:&XS�?��1�䕑{RR���mH�����rB���^4�����c�C�Ao>8,�;�0���I�GS����e�ԛ���X��"Kc`�ŠD�_X'��@�Tg߮�qg���`Ei�́��4�+^����s��A:bk�A�<C��4j8�[��K�N�3�����Q���?ym����<��f|9��C�����T=��⿙ jw�Չ��s4m�2�-�IF������خo�jz�]�G`�Q�Ą'`k��*(K��L�%��|ɆV���5!��u��KJ��e2@���P�Yנ�T{(����o1�r�B+����� ֊���Hڻ�2�K���*t�k��\��$ߗ���w�<DPK�<�4����#a4�i
�D���$�(��+�C)"� ǜ�K�\t*9F�=�Y�C>�B�G�[�`�7���7��{��!m� T.�</D�����=_�	>���@V��v"u'_�F�����-y���w�<���3�S���,6>6�Ўx��AQ<�Q����-JIN���3G}���8ѮD��@��u��XLC_9�W8�e!x�
@@o�l��4�C�T�*l�	��ST���W1X�|�ih���ѝ��qӹ��δ�P���	2��$"��[��T�3 ��:�JN�ȡ�ޑ��pD2���'@�YG��Z�L��4e�W='�sh6D'}�
qq6d�Qe���p�P@��3�U?��/"a�gM�d���O��3^��g���o��~���2��%)������$��
m�f�etFal�|J�!��YKU��ŝ�]\��L���-��8Ҁł�|6�8�z�D��(��!Y��Hk�nEL�,�h�L@=��\hr�5}{��*���_���8�|��q����9?JꊬVe��$�[Juǁ��W���r���Qq����_��|������³�ζ*��aU����A��-�l����:K4F�b��\M*srbR"+� C�"��s]���+���S�*�P���ׯဝ`��> rK.6�9�|��IAstT
!$�].��\�_��L*Mvz��9��.���Y�j_W%�V��z��ï������� �/�(�8b��p�Uc\��	_��ӦQ/�+�rYl���5�Z�㛁�9/�óe�4�lY����&����H�l�A~ڠ7�W�>��5C!�zh� KF<<�k���v�$��k��2�z�O����C!=�o8|�c�ͫd���zKa٬|[Te��W����Ju8����uF�Oh�B.���nbE?83p�M�H�����nF�lqf�ܼi$�:4�����?/}��&��
��"���9趘��q���G7��k��s��R7�p;�qO�Gc�^^� EɹiK�\s��@+�f���O/S��^f��M�Y�U�oM��V�>�� ��_H!�H�Ǳn!�b�f./�l��1��>]�b�HF=��oC���l�/���7C��~�VM,�K�>�:M��7`��	e�	��v[�� ؏��0��wa@5_�bN����\i����)�X�"�R�Q:^�{!�I��<V�FA���m�v�M� ��\�#�0��PJꒋ���B�C������M�c�h����^Pm�����q��`;i�����]ƴ��?�fj������{�=�{�����I䙶xb��S~�s֋2Q�d���)9���l�I�@%�DW��n�=`R�jl�F���?*RJ����3$�:[�CC,[�}M9��.��4��?�<�?]�_��7��i�#����b^�.ڗp?A�wD��}��m�Cd(_b�T�%^R-c��D zQ3�#�l�K�sB���}���F�|�	!���8������U�|x��!ߥK���d%!)�ũ���4��C�~�^��?E,9�.��F����z��u��?��g��Ȝ�� ��_�ڝfa?!���f�h�9��\5`n�B�q���)���Z����,$=��(�?��"V���F�e�,�݌�' �y��oR��nN��w7i��T��H[�ۥnqqqD��E�x��,6*�Qux���2\�u�k�RL$z��A-�Y2r�u�˷����M]
*F�ͧ�`�Yؓg=�'vd�r`��V������������e�{фTؗ��n[��W1��Ѵ�]�����r�匼�UD>�dN�T����`�&/�C��ˬ-s�ȼ��"G��-Ƣ���E�s�*f����O\�5H��K�OFn];રtA�֏
�W��$E���\�_�*6�+�9=����Ջ�A|_�<�}?{^�G�K�Am&����"����I�Eʳ֘f�=t)$�b�w��rt��k�����<�H����0�:[�����1��>Ԯ���^������O*dN)��y����՚R�߃���eU��V�c$�� գ�9H�U|G��褂��>ٝL_�R@��|e�L�~y�s_�6�}�--�_LZ�� l������ 'H�J'�N2E"��jY��m|��;h��.��Nޯ�-�0g��d�������S_�dM�xE��۱� �|\hg�[hlrs�)�x�:�|,���l�X_�T4���Jc :+���l��=6���[����3"Rڮv*i���'��1�p�)u��,K�B��bq��ݲ]����W;"�!~��ǃ�3Κ���R��H7���쾧�5�5�� X@�5`t�C?�k�􄅦�Z*&h6�L���꺩��Hm�|�q��qe~�L����M�U��@Iy&"+���p/NP���R4��G�Np����l<Z߉Wd���bO�[#�*���So��G�-@�_�j(vd:�h�]Ӑ8��~���|~���լ�4�#|=5Ov5<ݻ܋�_���"���3���5D~�nt��^R��ȼ�A=/P��/ה�!�.�z����a�r���eYM|J^o>��������G`�w�~�{JT�i��\�#��(�r?�ʢy�����P:g��?��h�Rx<!��b����s:3#'zK�S6ӺT�7~<���\��'���,��ٷ�[ĺ�t��@�1�`�5I�x�2~�3P��L�K��q��d�>���]y�Z���5��6�_.�`HS�������Cݗ�E7R�S%���^z���K�`�#����E��.�*G�Y7,�6f_eB(��������o�YQ����m^����k`aN*/�~�o�x��{�5���򋍡�
*4��[=��C��>�O!�.���A/]U�kl��h�����e�@_>w4ի�#_x���Y����PɔIjKXX���+�?�D�[Os���b�d����QF�-!��P"ɡY��Ҵ�.��.�Yp{�n4[ِv�l�^M�()�"ֳH��|Sy./����C}�R�^�H����{PI��ŵy��;I��rH,�͈��r=Q��_������=�U*��	����c�D�[
�ݴ3o�H+�w��$_�Q =U����j�A�G�֤�>?Yt��Rnj�	�-�q�SR2��Q�v  ���b.��n�ަR�^�#��s�+�_L��Y�xf�&G�#T0K���rX�L�-����J���MV��x���]�@�(��5��:�h�[轍u�y�+lD��憒����"�)~�a�s�ݞ�� e�CA�<�eW	#'_��܍����B��J<r���C�N�5+eE<�E�Ҵ�E����cS�`0ze�Tt�������@�6�/�zs�3�+�V���jY⼣�VdX�m�o�٢�0=��.���/�gɮP�t�羄��4�º0�<Q����^Ss�W�
K&w�:����k��IG��o��>�0���י�k�5zR�Q�G�#��[Q����]�0\���h�ڣ��e�MBa���N|=r;��E��d|��'G���;��Ɣ��_��n�5f�a�e�ɢ� �������Ɔd����fL:H*�M��p=c���:+Gˠ�K&j����� 7�	}��7�gs}͍tp�	ʒ�^}��%Н~�V���*Y6�0Q�M��bn��UF�A�X���8�����f�1��y��(U\��}/�b[�WŠ���^�A��D��[b۽��� �#�l���|�J<7;�:	�|+�o���<~�Ѩ�"O���E��?IN�Š���_��x��7�=1���ո�"?��Hj�� �n��W#r�&ux�\'r��|���DM�PL1��M�,��>�|S)SO�@�~� �~��>���k��b�V	����ge���	4� �Pw"RY,�^�l�x��Ǥ;�W��K�۶�tl۶mg�vǶ�ctl�c�۞ss_��Z���/;�%J �L'��_}0@_�L��լ��i��� ���I������VX��~�L�B%/��-m��m�V�蠻�A���>��3����'�T"L�0d.�;��	.��"��qH�hy��@nwM1A+�9�J�ǚ�ϲM�Ԙ�m�jRh�=�Dr#&(ʛǛfׁDz*�.�\�� ٞv��p>�nn�P���������m���G��"�j������7h�%����p]���)��'��|%���N���G%�6��r��e�(mgYt7���k%��Yt	�R�em��ĞYB��?Op�Ç�f��lN����m�1�#�'��ǷU�8�e,S� �A:��yG]$��m�Ir��a9�_�;ȗ��<T��ƕ�VVsٍ��d�Sd0L\#�>H%F#ċ��Wt��'�����W��Ǆ�6h4-���A|$c��b!�+�Mo���]X�,�u�z�꽺�� � �����N�xp�����	<P��k-,��y�� 6+O�Y+u�oV|*ښ6��I�%���'ЫwT���^R"5C^��󧊕��a��u:�5�to
�"of}�PZ7l�.���U�Z�*  �G���^&z�
�#ou}�2Y5	p�v=�1��З1]n1�ڐ�cz?�s�G�nw�>��1�/�Cmt�$�c��$J�*W�#��ê���3��Qq���#$���� {z N�� ^��'ր�K#L�ÛHs�2� |��7��]�E�0fz�Y�!e�~���������PpO� b�̙޿%���M�����M��6�Y��ﹿ�:�^<ij��TL��lQ)��X29�x���S]�2	�{I<��%���ٮ�C~*�]S���Z����C�m$!a}���R%8\�(�j�c �e�e�*,��� iX8���-�y�*��.��h�@�W��Q��L��gQ�(��NV���8Wvȫ�l*V<����2,z�g���B]ڤ^��$�-`�7��U��i�����֬v��5(
eM�,5��O C���Xo��/d�B�S�p��r��������5�عZoY�$p�/��?�3������l�$8țQ�mV����ؤ�*����Exp}-L������8�p�@h�a!9���y��{�Sr?In�`UA�ZLߔ�M����*e���,��D>�,�*'F�D��K��	΢�����o�q�Z��SC��|�f� ;�U[�JcN��S���Mឣ-���B��Yފh�*o�A��G�)�_��Q2U��Ɇ����G�<l C������8#Piv���!q)�ܑ���|
�����t�Q7~�>�>�!�aA7_6�@�:��2��8�5��S��������un��Cum)����A������M�U���!��WNIiM�/�OY̖��Щߎ8���h��q�c?<nUG��8'I5d�Xp��s���s����^�����>��8!朞���7Iv�M��8��V^�ʉ5�B>(#x�![�CQX8\�{����)�x�4@k�_>u�e�||B�����.p��'^n$��[�|4ۇ�*�pr�(W��G`�vu�?�	�������9�G]�[�D(�S!���9�x� �2���N-�
��w��:�&�Or�k�b��)֣�o�a+ r�mQ�t(B�a�k��,���6���0�0ht����@�c��K���ߩ�|��	������S,9�.#�Y74E$��ȴAUרMxU�����pˎ���V�g� sn?)���[�!;�I1"X�/ʑ!Ũ(w��əz[A9ѥ�T�A1�C�j����,u��yE�=Gl[�V]�t���j+N?�ht.���i[띢�"y�v�5e�t��������G��v�	��DDﮖ��fͺ0լ��&����z����1�y��q������w����1����3!p+m4�c���x/���X�f5�d] �=��I���<@Y�W�O�����ϧ��A���+��0�9����Z��zA��z�J� C,������k{t�m���V�bv��:���{h�:pe����'d��5����b����>2�2{@\�L=�],�6ԍt�]�T���2��u�*`R���ܱ���>��Px���?�y�f��f�Xe��g���郋��5�-���ҧsZ�H�E��N��AHw-9� K�Uh�H���&Em�d�q�y�c`��9MW ?{ gX� j<������4[7�Az���x�<U-�Y�5��]���u7J�]����s[bu���q���[L.��E��P0,�����𙰼1��0$�����
KW��, l�쎴�_=�F%��=K	��?n�_������,YdFD�N��^��6��
�>ZN���7k�NH�!��dVA��V��"q���7��m��F\.=�Yb�I�a���@[	�$f�@�����1���mߞ_�[fX8��ͻ���w7��~v� ��fMr\���U/Q8��q��d�c�) ��������iZ��}I+��9��D,ZP#[}��,���X+:�c#B>:[8�iC��ڦ����c(})�V�{�4�*���~�~YG�@��u�\����s�d6��� ���0x�	]��ڒ�ttuZz��=c�$ǴwJ��+�x��~��8ve��9�����D�|�1��5����Ž� ���LlU�0#h��Yuj�e��F���E�ȡ\��f��[�IX��w2̱ˠC�k?@�t�Ū��ڂvk�(�c�݉O�\�t�C�3y͔t��	�R!���F���ƭV#\�)ǆ�&�G0��������0M2�hkپ�>��݊2���`�TC���w��߶��R$������	�­
�f]��w0�9��JYuωo�͝��ͺ�� �w"!�Y��ĥc��{��f|�F��e�k���£Ða���ϐt���fީ?8� q��g��&OmI|���~�%�c��������a�����+�1Λǀ��[a���x?�X�?�B�J-S�i�#���"�.���#{�ѥ�n����o���u&�RdvZ�B���zY-���c_�7!��_����Q�81���p"v��(�aINU�l�7"�)u�mtY�B�����c������?��C��$3�M���g���I(��U��%��� o�����~���G���?�p�=S�|�A��ֈj�d��O���J⹧�)����u��Z�(���]a�*O"�]�/Z���梨@��ٻ<������T�-,^,�'Sw.���]��]�1������&��ݫmC-����{jW����n9���z�z���U�H���KsR�c�ߌ [����Z��+���p���;&+V���u���o�]7/L7o�h�	6L��_�}͹��(!\����԰�&�P���Y�|;�9�F���l�%��h�5z�����Z:��j�B;U��cd`Y���|�)�x-�Z�"�2h{��:P&�sٯ*���28�O�q���Z�����x��_�n�����C�s�؝2%��d`\���6��� __����Q{{$v~t���=�?@A�0|F� ~*EQY����?LF���/��=�63����&�K.�Ȗ�_�S���0�'�ѧV��0����5��ڔ:��3�!��]������^���1pE^���H.�ݸJ������>����2�wzb��y��Ú4Wm��<��ku�1x�׺:�{{��F��#$���7hV�11��� ��2uk��6�ظ��+w�t����]ך&�L(������I��c�C��@ע;�ԉP|ľ8E���V}"L�e��g��%"����KJ^Lo1*a���L�J�v8qo���<�t��{�q�0n�m)M�.��9h���Z{+����� �sc���&P`���F��C� ���h>��'��{��˶u�aӱbyZM���)-��`r`A+����|*W$�:�$��&�v%��tm��y�"U�d���%��
��C����7ZL�rG~~?<gd����q�\/�u���m��˪9H��uj�Y=�����J,�9�c��ܔ�ϧ:H��o��E�s��Φ��Ǒ� �t�����}R�s<�W�6��t��a�kH�b5ܚv�3��A[b%3&9Zj.B����D�������t+�ev+R��1N?P*��e�UUܫU-`҈S���M����Ma�(�#��IHP�%vy(�w� �=�8��pp��|���{;.�6����3�Ᏽsl�b3-E�,e]ƺ{_�	'�1PO7�s���=��ga��M;Nvs�(��Wi��r>]�P���p1#���S�n<�31i�v�[�8�0���Y~����)q�Xfy{�O��`^��@��#��x�ws���C��~�,|�G~ҁ�mש39���]0��oAO L�*��7�˚�e�,gpl�ͷ���T�碮H��,W��e�\�S�S�7E�	�H�ǩ*"l���;[��x���GP������cY[B�op�z<T��h���x3�)s�f�K����+����n%�>�x@h����������(`����'�s�����p=	�����yh��{e=���9��﻾JR�v*��dr��[[,lr�ϲ*���U��ފ�U^.�z!�u�Aw�_�擉��:��sP�Pȁ�6`ʖ����H�K�˅��/���
=�D��~8���HsE+�]��΀&�1:��9	��Ad	��fT� l��D�I��8�N���L���K4��}V�x��z�x�?�f��_�g���e3��Z��,[�@�>�)K��"��"�9�f/V�(<+��)�6��"�X��PE{H�;2�=\n�A]@���ܮ�z�#{ʲ�o��Ðs�,�:��1�@c	f�T,�*xf�tq �x�lR��/����M��z�C���t�Lsi6�\�������4V����j�r2�)R��ֳ^K:�n�uD�m��V�E(d�G���%:� �x 0Ԩ�
6}E9'J��[3U7��/�^O�/���g؏ ��Ia�ʒȡ���(�,�.r�J.L�j�A|��a Kv��p����)���h6�,�t^��0_G�X	�����&|r!ؖ�Y��N�j'���e*S�P,��`t.�<Q$�[�yQ>�����T�"�^��mZ(j�{�K�5Ϥq$'l���B�4Nloۻ;�EW�UE�kdV�8�Ց�
��i`�b�F��C�p�v���� ��R����v�P����0�O<1��y��`�R�3�zY�&uQob��)ܬ	\k}��v%p�m��8o"�V�1�Dś'�C��{���k�{�p�����^���:�+�TW��������?
wb@�������y��f�]�ϸb�FZ�������Fu'i�%kKK(�B:��k7P�C��^���(�-ۿOZ\(ؑ�s�L���&C5�iF�S���'�ҹW4C$�C&�Uk�t������'�O�5�S|{o��#Hڟ�h�3�@��?� �~<b�ە�Z�����a�j\/ ���9{(�ӹ=���i�S�2|�s�������i��0�==$*��U�+;�>~r��3��ܳز�wq�?/�C9�"y�!@��I����M�d���c��K4v�7��t�m�pF����{��<Ƅ7Pm;��S��.)ZE�4�Nz����D��~F����<��yx��V��@�A�����6[ѩ��l�/]^8����okd6�`��t���D�eU�Jq��P2,&�Q�A���6+1Y	X���E��h�h]MSI�l��5��n�.}�֖ΐ�o86rd(iC'��|�N�O�F�Bpn�O��혋�:��TQ����Xg�?$�~�9HȞ��e�Fl6���y:��K<��g�g@݈׊������L���fA��ꂻUc��sn�;(�ͼ�s�+z��7Q� o۹��Tj"��&F\W��O��a��R12Z*����H�O[Bw��5��"v^����E��v2���!&�EA�]�;5qdS17�p����ϔfg`�D�9�Y�i�+�/������h!�S��r ���2eb�J�f��P*KD�a��m^.p�*����,eu�,���C'l��Ŧ��zS쁛��� ݨ4��h���&A"��V��&+
�8�(�n(��c��ق��g�a�"$��|f� �����_t�bS��]M:���@�XJ�jF
4�*���F6{�L�P�ۏ�#c��v=�]���@����rɷt��t%��� Ʉ��:��s�G�S-O�p�v���#�D��ESG��F��q�-��Ԛ@b~��H<�' 4Ƀ=�I .ņ���X��!	�#�D�pS�T1��\��%D�몕��m�kxN;�X��;�x�Ӓ^�8�!U�e5�~�����n�����~z&h�0eW���б�s�ml��Q�D1&P7�������270ǻ��`��5�Ǹ��"��=RW������@O�=�j�����p9���l� �~���z�V���(XQai��wuu����	Qh��Vbks7I��(�����%A�-�����͆��M�m-?ƒ%lWY���\��\�5�;�i�A�c��/	�/
&�:>7 ���ԢA�X�X�F�����Ŵ�<C����7�$�}�51����Oы�#�M�l�:VG2h�Up��#奖 G,q.ӟ
鱟f	���>m���5��*O�`��3�aS�䠫R�:�d4���R�2�%Y�L�`�x��ռ
�h��~0Yh[�A��ª
ڳ�^��s��4��|#�PIO���u����4�h����b0*�\ܿEkۯ}ޏ�}!U�՘�g>�����ɲG2��K�`s������*�m)w�ӮuD�1~�U��P��# ���@�U#9��x�?�����1i�:�ߎv�qR�^�'hp�5��p�׏�D��4%r�h>3��m��fJa���80,̨Z6���:�%����%�^��Q�����;��������
>	{�g X݅�uL��,���ҊSk=���ƶ'��8�b�����۵/�U�1y ���ы��wk�6���2��(x�� ��Zu�`֊.�P�s�FU��N�/����2o`�OU�v�1w�֫.���z+��Kٸc8��n�WA����z/4���ѠmR���u��כ0��,�����`�׽�-�s��)��X����]ܮ�ډL=ҹC�VJy&{��`����EuQ��c�bO��w���@F�a=D�U{ʃf�0���������%����gh�v\��[�.�Z���>�9dԉW`� o9���dܡ��8J �Q�i;-��b�������s[9$�#�<���4z���~�e��&_�@��K�(y� 2|Q�%�ᆢ�5*����fo�#}����ހ�����dP|�N���g�}~���zݏekEu��+���]8�xR���GԾT�W�]ٻ���"�#���M^�tu�	*�Y��!%�wX?�E9��%1�k9�SÛS�W>�,��c����2�%]6��a���L�#c�����RLl	�+{Ń�9?s�.yJ8s���Ď�`�B�4�$"��g�f����=�V�VF���]b#�����!��^��P�p�qH�l��~s~|�J.�K��/ő�o���S+�ҹS����~G����7T��Ŝ�U���I�|���o#+Į�K��[����uO�;�_{��y3_>����HTa;�&\�	
�����b���C�5�Cׁ��ý��!z��?�<Ѵ/A��BA+	��B�|��_�U�<K���)����7%tu�.�����j��)�f�>��۷�A)[J9�s����R�`� 
�T���x>ɸ�q�y#9;k��q3����cL%����u�h#*���}/TE�������ZB��Lv������8x{����H\oAȇ��1������;qnH��"�2B V���q�Н�7�P}K��S���}�]x���Raӈ)�7�e�Â}V�X���M�;o�e{�%�0~����Dc���8����g��n����ܔ����x&���,�p>�t���0]�v���m'���@k�n��F[���A���&�|i0`9�w����4ʲV��k���A*
��GJ�4�^FZ0��uf:Ե)��_�m9>��R��
a�Br��x"��u��V���f�ù̅I1.�a�3k�V2��	�=n��Y��Zߘ*w�[V{t������ʃ���s�羀�v���L�}�H�r�\��x�x�.T�e�Ɍ˗��OIs���eI�/�7�D2�fyn?���o����R��{�`�	�l�3ן�����o�1؈K�k����rt�P���d	�~/�*��B*v����A=4+	Wm�Y�����Q����'�y�_p�P������ ���#��;��b=���_%Ğ��Xx�1���2[��=)0$Æ֤縡�Ɓ��y��.^�M-�(����h���LdyW�0�y�6/�a��n������O�MOa^-���/��f%��7;��y,��m�&�fRX�d-�x�y��E8> ��&sf��>��r�%�3��3Hu���M��je{��ʹ�����S����5ߔk�Վ�3{�a��͉kx����%���ST�^�X�ʙ�*���0�v�tH�X�N���L��Q�����Il5k$�#a���$ ��?�:�L�|?�W�wgnw;o��#%J$㍦��u�fz;$�^�*ew���Vj:���E�n�ݻn2-�/��L�P�O�vk�(�L�"�8Ӥ��>�#��L���o$�������#;�'�z�HqH&N �}b�u��r�os��nae�k.5a�)ծ��A��Dŵ�`f��Fֿr1��ZA2�뱢'� Qg%��-^�0L�+ot���+u���+q�G|���1��.��C�I����BAp�V^v��M�3�D�6�M�ɻ�)�U�����j���G�m%մP�O����F��p����=��S�d����՟>Nל����D2|��ު���1�R?�݇@�5��|`�{Tt���P<ciח���1����3�3D��Cх/gΐe�
�"d[��L�|j/�E������ll��z
M� �F���� ���EVtLO٘�C��+;�HW/݊hJX,߇?O(����B暋)�|�������E����`a;�R*	e��Qh�C Q��E���I��O�gr���{�����c�J��}|Nt����o_�I�#y1�~f]<j�c��� ���O����[�%�l��8��$r� f���z\��T�?H0k���)1�C�b����i9�lb!����(�h�D�W�#�ʽuj�U8Y+	EkӸ�̒'x� 0iN*�h��M��]�Az{�_[�+xV
Ŵ�w���p�bA����d��}<>Q�7�%t��F��YM:���EwD>��ߣ_eeU�볜b^�Zf�CA� �!p���Q#1f��($ȈQ#��1[4���$i��$�����)��dQ�c�ª���[A�k˳Q�յӫ�J\����gϙ�1�;�|�H���Cn��`0�P�ր��+��=8e�����觟���Xw����'א/g�!
���1�P��#^�$
���v��cnZ��l���!2�a���\&t��@@W���I�Y x-���m�1:E�Zl[�/���:u�de�~�Xb4ND�g~�m��5��6EOc>~��Q�0[� m0;ن�e�ߍ��?�&&�G����F��|*�=XN�?<����=�[c��
=�1ec,:�!_��v�}>IQ�2/�cgf�~��t��G�yT:��Lꒅ9G5���f�I��a���v�)%�h���G����lB1wk�t�x`0�]킲���D
u��d�D��(m�H�n�:f�9��W���2""1d��#jhR�����ӿ۝��*c�
F��!�-(�Ӧ�	s�懶�)@P]���<!���=W����GQCw�I�r�[�K���4.�
�*pCMns������:���Q[=}��T��}��ϓyhe���+g"+\��>*V"�����!<�@���l�3 ,t>H���p �c+c��ۨ�#�݆ʳ=F���*׮]�fI�_�>v+�Ȝͮ<�z��=�
�	}���"a4D$p�ś��@ղuj7���j�H��(=�qXί���O�j�wQAe�U��aƫS�%n�Ґ=E�\�s<�hl�4@��af+Ё���f�o��#�L�M��k~%�������g��W�Ti�g����T��+n*.�v�S��V���_�<ڢ�ٖ�zr���o�������ujV�:1�%$��a��$yb\5@���gj����%��΄Kֻ�hP���"R4��+3�45�}.�:�t,DZ`�T�v_"g':�E�G��Oq�D�('GR�;�s�F��օ����v�!b���'�lk�b�����  �/Ւr�Wv\���NoB?�x�m�c�/xS1� 5����GT�&2Y,3�5�$=�RKI5w�:�"��a`rŖL>��#�Ē��8VA���>0�N�'i�"ӕ�Kca(1P"��❪�/-"�#}���):��>��f2�I��Pi�_.���� �63��fF��[o���%ͮ5E�N��9��:NN��Ú��==���v��v�����y^��j���oc�t�	�g]e&�"E=�R��#|��]�V��>�7㖀��fY�=��hPC3+��Ֆ@צ{�#םO��ӂ�2p�����ɼ�飑9%�3��h}#��R^���J��fY��'~�B���Hn���/�Y�͖ÿnꪊBn���ח����l��reI֍x=��_�a�iu$�0��W����P�[#����V��;��IXfs��B�X��F�<��.�Pr��(Pe9��LM&���q�e��Em�����?�VZ%�C�T��
�vܔ(/����85�_�	��W0+�E���B c���L��^7�dB�(N�mJe.�P�`i����/�	_�J���7�Td�NT�Y[��Oc 2x�I�ys8P���>V��xW w�VC�GaxԠ@M��b��"��p�]A���{Gr���Yԗ4�ޏ,������Q���+�T>�1{/�a^���PY���p��bVm��E�0�d1nV;(g���h���nnΈ̆]���To���5�CP/w8W��F'eIDΥY��F=��
uɴ�aTO
�F�A�h�-�Zf���<�BT��0�^�ǚ9�B�3��+$��ޚ��1����������1B+S_�v��2�M�W;!bɤ#�P�|���
ǉ�G����y�S=�y�~�j6X�p%(�ˇ]a`@~2������1��ڧҬ���r=��[$m%�
�x=#gٰ�@�SG�2O��"Q�&L&��0m���#�S��Jn�~�i|���[OO�t�cT�/�	�܉Tpm�[-�=m�0ѝ����{6�(=��JEU3�rH�V�h&�_��*v�?��}?��2੶r0���LD��+r�>������+p�'%;�ńö��V+�L�^#���c-�ʩ A�W�*��ɿ�6Ub��>���.�aK�(�jOי��$G1
 p^|m��]H��IN�%�CП�����w�����@"�ڲ�)_�[W�@|��ə�d�>���j�����\���#�V�~�/�
S.4)^�AGN�����_��3@鋌�@/�)�l� �ci�RP�B��jZF�Xۥ�x��o&p�P
�t���iԌL��j���*au��,%���$x��C�v���k��j�0��+PpKULx������葴���_�`(M��nsB٨T��y.TV0p��U��)��C�gb����c������0�00{u���������f#<{��Pr����%� �`��{?X�������.Gܯ}����&G���_=����qY����ãt��H�֠��rI�-�s�QZt3V[�$��{�ƷJ�Z����?�����D#(Q����׬�)��c
� ���$�g�NO��1=��qDr)l��B�i�Ph.5Q�|�G��Y�p�e@�1"G� `�4�T��qv�������W
]mm�\��Բ_���1wlC��!�����B=����s��vU^�/�#���G!u��`i����Z����P��
9R6�:Df�����-�8ю�Sє�*~$k�e�
��r��VND���P;ɻ��-��М�d�7(����j���g>����o��uZ\�.�׏�MM�quM0���2]�5ǯ{E�5�{<��*�v� c5,LfT��� �k^�h���=�B�0�9uM� j�e����ńs�{{�EŬ�����K3aͲO�����~�s7�nܢ����\���<��;ˤzII���e�\4ɧK]@+����-L��-^*~s��r`�q5m`:�4^�#��ցhk�o;�q��{�v��K�]�=�2D9ʲ�T��m�N���J�CN�����.Q?C��ٝ,�E &T�*;�	�f�]Z(a�a�#k�l�>#Y�B���{���-�~�9�U����>sW$��^�yƗp���5dG4�Xۦ���u+���w�i�������	fG�����s�踻�ٍ#��A�5�W�=�~��}`��l�3;��X��a��l�~=�@���v7�z���·|G,�V���=d3��sf���F_I�|�9�ͥ�{�d�?6�[�^�dGӵ���GrM�H�o���Z�([(E���թG���f���P�Q>A��W�L��:.��M�Q���,%~����x�܎�O7([f����ޟq�|������u>Zݨ��x{�t���j��~�����d"�?94�iy��:x�/У;\1T�z,��݆:֬��[gݓ7�eg	R����Y�$�͇�c��׷ɇ�G�a��N#!�|�q��P�XPy~�Z^�L�,~��z�٪W��R�\��ȫ�o���pEz�̍:�V�
11���`%n��}~�f�^��%�[U0HN����Z7��p�:��߽��m����B�d�~��。s�6l�� !<f�1���w�|VoZ�+e:�{��X����R��8�-/Y��f��z���t`���E0�Xtc�W�W>��L��9�4�H�:�v-H$��)�XR[(�)���v(�<����} p�"t|�	K��}�� ��wN;3K���Y��u���s��l�bpI�|�������B���Y^k��a������w�/��� �¥x*$JNN��6PsP޷���k���u��E3����M/I���~���yո�dT ���N�ߗ��
����EK�E�=��ĳ1LBo��*rkJ�`������@r�_g�T�����!��6ڹ���qk1WL�Ȟ3k�jY�9��@��_��Z�\�CY�	����ச�`\{�y�p�kj�܏��y�9�C����s��Z�wa��lv45� K���Yr|��x�����
;��O��<��ԥ�vAo/ف6��~��U�^��qKŬ`��A�r���(/F)Sw�N����fǑ2O��b��� )��1�f7���`�'��q'Z��ɤ�]�chYF�XT��&�e3��)M-���w C�)6�h��ڔd�qe�����O8��0vewk���d��s�A�����ruk"��m��T�֐���uיf��危S7��� _����Z�NR�35�>���^sZ>d��!����P$.2չ[/�f�g��J�v�d�Y)�\���\�_����zk����}�ѓՃ44���߄_>���F�YD�⒉_m�	�]�a𬩈���%;�V�����z�D[�f�j�����t�)�J��M=�T$xX�D�H?@�"L�]�41��Heѵo����4�c��� a0���r�h���G$������0�̨��3�TߒD����.��j١�0�RԦo��G]ů�x�s��u�/ӈx'�ԗ�6&V�)Ȧ���U|k"����>� @6����c�nQ[E����1_� c-r�u��,ƒ0�^�;���K$�����e��+o�q� _����NE����9����%�=�C�������U5�W��)�l
��5	i��/u�S)߶P@e\c��!�b�p޽��Y��[Z�Ȩ�h�\슃�D.��{�"`7j4ai�»qo<�WS�����[*��;�b�T�U1����|{�m! �G�2�nW��cOmJ�k��'�Ծ��ַ��ғ��i�CF?���m�
��������$���#�YJv=�-1F��[<�"��CX���,9i���{�F�n��{"M��N�Ff�;H	����t2�_��r���8��檜|#���M)!������|�5z��tí���Z9�d7^���Ϻ�bD�y��CRj��]�G2�3�K��]�W��V�r��h�:n��~q3��+c�
��BؤQ�E�U��i4�k��w��R��^�W��cS�{.�&�O��$��ظ��E�����"�~�4�j��|H͔�M�<�h4Զc����v�ي��?��'��C���cf�N�D�-�e�
��ǁ�'6.N�����B�	�g&����O��D�wƟ������Cm�5=��ߑ13|HXv[q��
I��Y��u�x�|�~���T5h����Q�&�^V~�j5�\����w���.bf�{�FSO��T���{�R�ɞZLG8�'���0�Do�bC�����m-�g�y+��ϯ�/s���;D<:��y�ET�~�GI��l�3%޲�m �7S3�d܇.n �Z[�!b�[AL��-g�J��^f�$��m�i��!���{ը��c�5Ie��dN����	�I�Ӽl�9u"�4`�5�r��FG���:��2�����Q����PQuR]�eY�j��m���"	q�2lB�>d����e�U	��@�lE��	�4�vl��0N:�b�+T�V����ㄦib��ݬ�\�>�М0��J�9��7���r�-4"wxir`�i�~���\�ԩ���s�L�������M��/MB>K{���hR�$Ԯ��n-kó�ww�z���b�+Ү7�¤��&Z�wu����ɑW��ĎT�T^���UiK��?�rȁ�+�� y�UT��م���fAzt`���sN�7=����t�I���'�~wYp�H!��01�S[��>nb�m���T!�|H3�1J���$'���i����@�Rm3��Jߒ}���n�p����؆�Z�u��X/�h&J�#���FS��մ��KQ�GA��dB�e|�u��y���&������r4�%Ħnm`�͌�K�l��;+��T?�c�E"R����&{�nC�&^�]TF��6�`j�1�l����hs���*Y�,~
N��ȓ���QmBE#��3�Z�9�)�7<u�v�#Qд?j���̏��V�edbP�wZlȩ9��$����p�^PQ�'�����΢��ضylj�i�|+�n�pm�㎒��2C��Y ��-.v'* �ϴ���������3Q�W�z�Y�T,a�<�z+B���̣n$���l���1Ӹd�!���K��r��FS�2�0\�:�"9d|�����J�����F� �2$��!�d]���K.���9���Z�b`����e6��7�MhۆĪ� qFr��E!kg ��kK�q�js)9t�eqGJ�Re�8����`V�d��
�5�E���O�Mi9��W�A�	ۖ��A�����'){f_J�>�>��c�y1�fV�Y�q��N:2����W�KO(	�)OwFt^@�Y�����[B
T{��D���哛}�+�1����,mX׸�5�%$+Z6���x%���T�9�g�#K�����tC�UH&:w��º���T��~��W�R��H��z�i�7/O�bL��*Kq$�dt^�q#e�U:_<Av�O�^�"��)*�҆j����ݒl���@��ȧ/2�`t��y�-�920O��-��@�?I��-��W���b�����Zj���4A^��!�<岣�s��f�̯���E$f�q�̦� =���|�U*�~I��K�'��!Ġ���,��V�X�xهò%�ͱl����F�KKW�Ӓ+���(��buנ}A�[R;��p8Ͳ)8�&����hZ����Lv7fP�M����������V	�E�m�dO�m�dM��d۶�l���n�d�:5Y��������/�g�k����o�}7�<����Q*&Dٵ&J$ݴ��SL�!�0Gi���z?��4�3�r��2�Y-�� ���j[�r�z���;��L�8Q9C{���-���$��AF_�j�Gz�$l%|ط�+=8�p�Dǁ�[(�Q�)���_JS��z�q�����\56?�����VV|:����9݌�`�7�aV��O���M�"0�*�nO�0���Ј�3c���imVtvǗ@F� i	�=���Dji,X�Xa~�e�4����*�9�񶭶lH�`��z���du�Ҕ^�Y���Se%;B�-����\VV|)�n��/n5Yy������b�V�J��� d��o�F��h�:y��$

Z���9 �6�����b3���1_���VӹB��_�۽i�(�Nh�f*N�o�O>d�+�1��J�j�憓���[��GDq������ga���E� M2$��d��=A�Ư��;�n�hݰ_�9� ��\�~'Z2+��t#���H:ٮY��������=w��Ŏ+6�؟� ����/��ML���c�[k~JW��_z�]sX*��]Y`�ƅ�>I,�@o$Bc%�#��@�&$�l�M>��	��ZR����;�c*�HX�3C�O�|��S���,E�밖�	PM�T��ݳ�Ű8�r&X���S��n�ѻ��/KZ�]�i�]MU��$�Pzи�����Ca�A�}�BMi&&��H�2Yf��:�?h���v������ӼD�5�AD0r�rA.!ά�;��b�p��w��ڂ&�B�(��@e����k�,6���������e4~_�X��h��g�u�;�3(��k�:�R紹k��p)G�ų����/#P����t^��)��
��N��`��0<������#����Lo�l�I��lr�"[��M��v�$�=�o�/��&��v��6N������ę6��b.>���h���)&9�ܙ׺�������i˷��5��Ґ �fLޑi�`�q����ɂ�[�s�􉇄d�0 A�(#��b��M�^��t������TC�I�H��Z? B��-�V{C������k�-�bV)�1չ� ��-��!��k
s4��c7˰7v�Նv��q �������e:44��p0�X���j�cl\��Ƞ���GY�R�8����1n�ޭ]}x�������;�>s�;?�#y��Ep��$����F��Y�f��o��g�1Z��ct�UN5�=����\�ʆ/�(���'́�6��d�#�cCs<J�N+	�V���:P�/���02Ҩ��]H�^�O�߄n�_�;�z�{�C�������-+M�3	n�և�ǿ�jѾ3�����J\����G�y���]^Ws/����wj���R���� 6�0:{�c���gĲ��p@��!C�Xy]w{y����
��/��Ӧ��+��x�Ŗ-=m{WL|l���޴����^G����|������{I����݊�
�A��؇����Η����ޜ{��45 n�}!��E��� .�rn�1�rZ �?���֙�~�����u'*��>�ڑ�^����պ������q�'����Z��n���0x��F�aa���y�y��0>��3�sf��!<�M����q4G�/�X�=�]�&}�ؐ�,�@b�t	��d���k��.�B�1�l�d���F���|��m�@����c��~(��y�Qx���O��W��I��Ŷ�����+��vls�p��U�9��[ե�0t��@�|��+Y늙3���� M5��F����o��ss�Z��Y����Tml9+�~[�ܚ��ܮ��r���a�U��@�k3�h�~��H@��O�Ĺ���&��|j)��	��-,���n���P"x���D�Tn����H��r��7�%߽EO}3��f]D,K'
���'~`�.c?2K !K�#���=��%���:�i�����c���3���1KB��Y�po���u�F��!{���1�3)c��P�W���A��?���N�>S�&41�"��|����;w��M�XV�Y��i0��������n,��@�JkH�w�Z�;1��r�zR��2z-Nm���x������yj��Gu�H�VUL͚ɠ��~iW9-��F��ފ��Y}s����h�����p�Pң�ײKO|��0\@hTv[��w����5�^����!�s�����c���d}����a�u��=)p�뵬����
�K��Y2o�!O��"���|��7ע�h�V�z�x2�����"�&X�</��T�:��q�*�-qʹ�Y�ʅ��%���c�|Hh�,��в������ן�Sx	dCrl��gY.�5�2]sw:"^�	��1O���6:���+}O=`�y�G"��j0U*�����Fj�M|��6�߰s]��u�F\]�>�c�t� Vx���N��R�ƭi��@�����'�a�-��6U� T�)i�r%�%�~�6D��j�ǯ�F�EWBC�5���W�o�ˈ���ׇͧ,�C�B�l%�눋��!	���E���x��}��yKO����$y2%�K���w�c��J�}���:�Y$���	;�Pg�Om`,$J\�4.�on?|�T0G^����)[v� �F%oEz	�l�#"��g5�!� Z��ߐ(Gps�ke���A��f����s`j�!R��=�C�Y�f,�����'"�4�Dnd�z��5�nR[Y���0$�c/�Ն����O�̎F�Vs����~8�i�M�v�l��"q�5����Ie��i":��͔�J����c|��IM[]�5��u��oMu�+(����]�ev�\��t��C��M X]�؋k�\��MA��%��v@C�ͮkW>�In��MJi#N�frϑ}_0����\�&Dя.��͗]a���q~�/6Ex�|c�>ʙ�\s�*`����_��`�*_����E�d�H<x�5 ����?��i��q�n��8�V�?��'~��Md|Y�c ��̴.]
g�gRN�?��Q�d�I����^�������ZHr��0�HEb�f6$�4�X�L�M!�+#4�>����DÓ��]��)z]*w�w���8�<�&���~��{�:�0�$��G��ҧ�S��	�o+\�I�HTb������pӽ�[5q\`γ���zb��Ń��ϰ��z�ţ�>� _:�����*�sy�n��ñJ���o�2�<��H�=��g`�[:OSSRƷ	<��DDoHZ�+Ë�xqh�l}2����H���H5�v��+���_�e�o~x��J@�9Q:Ziٺbn���r�?I�l.�e^��9���d��ި�뉅�����W�Ѽ�o��4(�cL�e)����CQKv(��:z,YFL�Xj'�6\ۉE�6>y^x�7,�_2e�t����KZ���R^�|���{M���ިT0f��J��:�O�^B��������?�O�'p�]�J�ۑ�G��0�^�U�Ο&~x�3����D���_�l�І�J�FV�!�Qe��^����&�IJ��L�6</U�����lw����*�0�\�(X}�w��~ש�����ǞG_D�9H��g�0�
1�o)r���s��.c	?(k3�!��6!����5�,�\�j�z~��tjU�$�)������ڟ��y�^3d"���W���Gh�B��̠d���"��(j+4��c)�&b=���=��w^��Z-%c���y|/���g&�Wϻ�����[}�B��x��������+��/\�7��S#$
M���c8������*��Iqd=�xB^33llB��:���{��wPJj�HXe"�7k}��*��@5�S���c����!>�Q]dA>����I�B���N_�-P�";l�P�eH�TK��X���hg���;��p�}��4Hak��2!�������mzy#�0��.�BY[^6�o)��Tt�����SEx*�?���@�?%~��sK ��"����,Yb��ӓ̜Q�ê�������&�l��@-x�6����wr۸tbp��Ի��Hm��9���]|$�
���bS-Ap���h��I��R��=m��:��l����~�^��f���),�w�O;>���J��Rϸ��~��	�(���S/~��J�$��i�Q,�q��7����*�~�/^f*I"<�*�D�t��'�L����3�`��&�z��w���*�+���Z!�i�"��ߴ�Jv���r%���0���/^�| �z���2�:��Y^l���W��IW�jit2�X�����N���77�KE�����F�z�� �'U�
%���kz\�4��V��xu��l���g�v	�`r�נ��db �hHHL�����L����=o�#�<��?Vw*���{�D�������|��%b��\�T��=�i��%��"����Y��Y�����|��i� �?�2�t&���=�<�2M�o��Y|�ގ4÷��ߔO�%C�2�M41:A^5a�m{�#���W.;�e�"JX�Q�b��؀R�B^�1u~_��+2P��gF�x�P��LM�����(�X�C:����M
���&ȇd�gU"�/�n��*����q��m뗷���ɤK�CKQz�Z�nv0.��N��KX��;�ZEz�J%�K�l�O۷W8�;���y��B�j�|��%*�SM���5o��9���X,��c؝'��x�ymQ��n3�ӊ�`�1�4h�
=Œ�\����7�� J�r%�]0�#8 %�:)ܜ����=�א4aY�V�8i��Tq}gߌH-E���<��d{�;�9s���Z���~>a��>��g����k�	���J<�i���^� D��v��6dK[gԗ�cJ������5�	]>��5t$4�rn� ��O�<��h��>�q�h[�T��$��������I�$���M(<��Е�I-7��Ĵ��؈)����V���u8��bFD�݇$eX���3�j ��������ŏ4��xyy�M��.��c����Q���%��q+#ہ�2Μ��� ����lM��"݊�"��$���ݛcN�����9���	�y�L��Q��.O[2|I��RU=ͬ)Y��MJ7^Nҡ��yw/�J��4�Y���s1_��%�ȶ"�>��*2̼�辌��j��T4m�!4�
��O|j
��8�yJe��z]
��[g�ny�e��YK:V�-0o����r�
�u�ôS�O;[��U��w�a��7��p�q;P[�h9��cH�~)d�ώ@��	�⁢2P�W�u���?�c�j�u/�g�	�Kvi0,9��5�� I��xy�7 4N�Adj�b�{\s�i��Kp��?*Ys%���gr�ʗ�d �ꘋ�@SԈ/�������"�7<�>�tu_W"��aC��~�O�f0��G�x�>�/e482���W���zR%sR1����!��:�1��H7h�+-�]��1�j�W̒�K��G�4*�h;Ւ���m�ץ�E��.���態v�˙Ҹ�0�`�����l�N�MzT�I}i�z��0�\��m�#��b�yc:���@��u�U�f���P��7$((N5���ע����lR\lTyN��Iz��I�1��Z=��,���Zl�7�6�Du�;ol�E��9�̷�%J��o�>2p�P�\h��ژ����C\�[���M�v��G�_c@
�u��,+��X���D�料K��,ӹ$	3\�&J�`
�[h�Y�娜�a�p�t'f��u�4�^�]-��T=�z�$���ѹ�OlJ������z5o��)P��x���_֬�钮��G3�6hGVƮ�̈a����������z-���R����,8��������'l�5I˻��	ߒ�ˡ��r�`R���@�3,fyiɧ��܁*�mP�"u��H��}����-x�/Exah|�=I��!Mo����ml���� ϖG&�؛��N�ޗ����� FVU&K|@7 ��t��n$���rd�D��56ɨ�����~�J�n����Y��R���Vgq�+WS[�t:�
�&z�֬L_�	��$�{3��?�jaQV7�B���D�g�̾�
϶I	7��ѐ��g�Y�'��o�>?W�3Y�f��-34��`p�[����S����RK��yi���e�A����ȕ��mD�������?����'#**x�@޲�� ]�_9�_{��6��<�tzP�?OO{�8M�Q�%���P4�z��4�ZS����	*=�pY	~iVb�n�4j�pʍ.��%�"��.�zTD����>�	�¾j�=�1�-Q��s��S�]�<�a��E4XN�!{��h�Dk�#"��7�_��ĺ���Q���hbĺ�WCb�Ŵ��ۋ�b%폭<��Y�j^�3��0Թ�s]�r�h]ҴU�ϠsW9Z�UW�_�J���"oZ�x���#|�do)n6֋�X�LCx������G�3�EeXN�=�D�����7"k���Ai��%Zt^��>4����n���Re=}*\]��(��Py	�^�ը�e��&m�-�ʎ1̥$�����N |������u���1A��3�6B�c�^ots�#�4/��uE�$�~&O�L(hE�Mqh�@��~f�B�K���Q��/~d�_�"��&��_Q���ԒyL˛W}Gbo�����<Q�o\h���c����{&��K�Q���"p�d{/\r?�u 6�v�#�O{�s�^}'���W�U��,w\�����֟�������^�e�z��?N
�zW����nM-�~^��?��r]��I׫c�.	O]W�W7���ge�@��%����?�w���h�|X5����d�dŤ~��V7b�po��<w���Y�)��QA�)���A.R�Xn�;��m��-;6m(��{e�s��"T�bD�Y�8 ��Y �y��H��ue؎��=-M�Z�_��g����*�2��>f'�ۦdg���\�����6jf���i�"�G���ʀ��a��tI~��S�X�|��뮐���H�'������}I.�Pc��l@2��{V֕"x14(F������^����|��C��,R�
�_L^��E����w;X���g���r�5��S;w�A�Imx��ΐ�ï�2׽�?�T%p�[@�0\�9���rpO�n�����W7���i���}��1i��6�h�4�׾k"���Y��`;��
�!�{�׭D���.��_Z3wi��8f��b���X~�Qbv$!��.��!�jZ������N~M���*�׆����[����629�G( ���!h�4���\�G�y���9��=LM�f(`�r��~3i2Ȥ���s�A�8�8{a̙�<[��32^F���V��o��~��/E���l?a��m��w�Jӆ���<�4�l�}����ˎm��y7'���|m�M�y������:c���"��1��Sym޾����D=�f������ݜ�e��	g�i��6i2�/�������ƹ�ވ>���*���4	�zPr�
V斓�F:!��nQ�Y����}q���!(A
��0`S!ɴ�������P�U�h�m��4�tk���O���T���m�9�O^�?쌡Q�H�V��B�3��f��:n��}a����z���<8��1�?=���W�?+��kr~6���������S���i���Hя>��=�z?�:��k���©�@cwm����t���p����
0���jA��":���G��^�����^r����s��������l_t��'�+#�d cC�:�V��+̝�g��������(� �<ɍ�{��Y��[�;q�xN��0��J6J-F������\y�B}\�|>jS[���7�������O������������.gj����G�_I~$G:�7��Q�Y������'�Z��kP��W����Q�n�zm�����"ev0��+u'�=JgOv&�2�IY��բ�63B��|��^/]u��"�+6"�A���r�:�X�E��鳭~ ��3k����z��r�~.�I�����1�`�y�t����-��4�~�%?ً�(�l�y�"��&ͥ͸�3�װo�4�i���HYپ��$�ж�A|���C�]]wW����
}�1O��:/u�G���is
� �x�8!0��E���iۃ<spZu7��:�.�"�x�@���U�_z���L���Ev ��k��ȓ��ѓHT�{dҗ�k]@�qO�	��6�N�	y�o��z��"��e�����5�YtJ0,��������N�R�]���sfx���F��\�o�\DQ#�U��h�"�t�~�3}�ArURgn�?��JrDS�����{��rț�`8�J9�+�@^�9tzn[��u���G150w���j��M�W1���iV�!��8u,���~_P�Z"�A�2EՈZ���b�C�$�R/��h��ܮFg�Oj3Ә�nz�0��0Ҽi�XM�� d¹ᒼ�"Q�L �����Kڐ���s�,|�@qi�K�qGWȃ�a5�!�w�����/���=iE�s'���В`�:�?���5q�|��83y�GEs�o�R�\��Ȩ}��� j�5�{�J��:�:�q+J�"0���ct�\s�ϐ F��p��=����k�,D�M?<aC��1����kc���k�$Z�;[Xa~��"$M��V��<
�gT~��w����	iO��^���sN�Rn}�tf1�"�%
G�ÎVZ�cr�O��m��9�����>?z\l���
9|�HPpK������Rj�P ?��(E.��h5h��0��0�1�1��Y�x0�}Xԛ��x��p��6�L.�g�mqR+���~�)�C6�����[W{�$֦A'��#�2��lܮH��ף��K+f!�	9�A������b�E�B��Ċ�Q�3s�>.�L��΄�F�J�s�j�B����0�� r�pÈ�5�y��k��5X�4m�	��� �-�ٟ�Qm�٤^�܍Lk�. �w���z��Z�˚���1�X��u!�aӡ��x �O'� q�(Wv�p	0=˫��^^B�����L�q�фB�&��V�0���w<�2�"fm	#��^'W�dYy��NW�?M�R-�/شu��$/�hK�&l()T�[�E���aשְ$�T���T0�C�ǝX�f[(t�� 'q9LE�n�����ͩ���J|v��Z{��+?v�\ �F�Gx�	>#'|n�Ӓ���Q/	��FV\?3�RY�	�����{�M(����[(nj]�v��!�\�/���"Z�
��ufF��^g�	��J�(F�G�p�E��I����#8�����SG��fx����!�Ҳ����"�4�2�����C�� �N'V����V\z�quX�8����tP�f5��^4��$W��� �.?���f���U���N���/���u�� �=B�=�]e��vE<9&�J/:DEG\E"�����?j)���.��^���EWޠ�ģ�,!��#��׮��i��"���"*R��������R�c�3�����jU5�ߺ�'��� E#��#a���J^o�����䨑`(	(�r��KjE�gZ��=��bV�q̎;�<�N�#ߘ�<�1���\m���A��H+��:��B���v����hZ�`��`��c�
p��U-�"E��� G�K�cݟ")�dRh����a�,�Ȓ��eĠLarL�C%��1�W�����y(�E�s�!Dy�!C��a�K��'��1��q�i��:]� �cUn�q�މ�l4?4���#X��4���5���F�2���k�I�,�}�>�·��9�22U��$i��GzD��Z,�=�1�!u���$s�9:�8�ɴ<2wk�6A~�.���g����]��h-�(��L%R�l�6xwɲ|�m��� ��}��)j���t�_jf��:��iB���������Jza	-�8:-����Ky��j����G,.A��JQ�2-p���2�<��@u���%� ;z]�H�_AL3�a�����o$���V�/��d��*�P�������2鼌g�F�'�:��^�/���^���e[2�҃v.n�K^����|��p���\lAXL����k�R�v�� &�F�4Ȑ�X~�f�̫"uH����_Y(�L�������$�?t*�BԞr�6IO}�/����uz'�*��_���R�Q�o��8�����ӪM���uM}R���~��qŐ*�S�?�����f�E�����.�m8T��O|*��OK2E�zz��ǆ��Y�5�:.��E�Q���ˬM<H~H��VҰ0}������-�J%Ag)��=W�2��{�O�~Z�����%���֙噏�2���Cɾ��]V>��� ��w{-�LDD��
�3�7[[�Ps�skE�I`W�/0N�1��xZ�n��%��q)��/a-�Q��[�D��OPGm����jO�A�G�e/�6���'��U�n�f$�#��b���AOr��G�s�Sj�s�L'���Hf���� K�g�K�>jX6�\;ZVX	W��y��������֮
��	5z>6�@@&Lz%{��M�PD����U6�]��Dh�8���VA�4��HE�ji���[��u��8KG�yJK�̤K5���[A^����#�EҸ]�l���H2�e�F�U���e�{\�%�� ��M���1#�Dĺ�"ܵ�Oq�G����X_K�{��`�7�T5���������y�4Fr��Y������ā7�g$"3����?ߌ��5�C�e�u��?�U(�F�Mo�>�@�M��&iۚ��ȑ��V�K�l��V�cF�h��eG�������\���<*#��8�s��C��7�N�
AK)H��у���U�U��λ�@�9�<E�8vD:[����%w�H$Z���<�Z�|5��F����,��R`�L֙��Jso[HZ�%�0�Z�D��������7�6��b |d$�`_ԟ7�_?�
'�X�&�f""�fWV*{@�zr,��Ӫ����?�؂$#ъ4��'G��Gɴ�6̼�ʣҩ�j߲ �����w����3ӯ�ޞLY�n�Qu����]Ĩ�|@:,�h�����F�]7'%�LE$ y_���j�45���.�i�0S�!(�e���j.�R-��w9"��n�����vY����&[z��N��4���0�~!������" ����` �f���G�ql�`�
j�`����?\ ���~y`���Ъ=���h��m~�1$[�B���V��ss��c��"�����RƝI�:F�V�;���g�xj�82#oo8MA3���=UO��S����5��"�&v�3Cڅ�1)K���f�K_�2;*�M����:{�+j�AS�a��̺�Ƌ�G#�.NBxu�V�u[��������w_��b}KԌ�9&!nn�:E)��.o@p��Â�Up�A�yV�1���:Z�-U2�.�b1��G���=`(��3�GD�k���#�5�XFh��´���� *k�?6����v1p��#����yJvI��1���Ĕ�\��F�2��$�t�L��n(�SL;�8A3;>d����GG�,_Ҭj(GY���c����G��"��L��2Y��q�):`7xu	��a�M�L�ߩ��-�KW)�f~WFz���L��2N��&���������?�DfL���K�*`NkibF��t��a����#��*��+�h���-�����0�[�׿K�e�7h��
�U,�0oI�G�8��Ү�wԜK�dN��e��!vd�_#L[�Q�{xz�k���ۨ�?a�K�4���E0[6����VUY9�`�2g~[P�U�6��� o
������j�*�� y��1�mf�jb(��/ɕW�ZJV�V�ڡ~.IZ��|}3Y�-
�cݠ����,���Q�t���3��{os3�P�3�V�D�v�s�]c�%MX�.��%G|��y^Ɖ��6��ԡnT��`)3����*>���:�ԋ�*M{����[&?n;�>�������3��F:t�2x�����"���2�_�ő4mUc�%�]��G�&G�f읮��ֹ���z�٘��'����á�B1X��rZ��]�F~9�!8:��p�=�Aߍ\�L�J���7�˕;@[�P�v�5�Y���:|H���gg��l�����Ź�۩�_ ����	;M
�I|�P���O��
~�\��W�?�[[WW7-��j�֬&��&&qh�z��CRWM�Z7�ot@|�6��5�ҼJ:C���XF�跍�1�s�O���nE~��q �Ar�/�[�~����������$Eq���3{��z\�.�tڗ�tP$��^+��9J9B�r�$��� Q����0�Ći�|�,Ί��#o&���@�7�
��N�40�%L� xX�֔�}�&S31�''͜��S�\pn�ABS��CC�T�!VM�ͭd�}a7$
�ͅG?���n��~k�u�"��yB>��E}�����8`�S�r��A�������`� ���N��-36��Ɵt�\���_�ו@���(��e�7nx-�������7t��t�֡�m�S�H�vJ�x�a���𬿆�i�-xD�+�W�2%�{�0�0k��O�+��"\�����P��@=ZH�`p��:j�΀O�*JӜӦ���������-��tqp���9��&�ۨQŇe�*��f2F�ME�[����܅�y��w��0%	��j���F�������Kw�>pq6$yy���R��#Dʦ3C�/�cx(�<�+[��t�b��F��b��Ъ��K�RY�b��l�1���wUӕ�^�	j�q�hm�����P�3Qk�ު��;��p���I0�W{�]�bj鍊~�$uF?�k��ڶ��R�	�������9��P��$�����ϼ|�\qLر�-N��b��_X��-S�}��Ok�;�#�c�3�����4�4̿T]8��8���H��v86�{�3��U��KF�Sɫd�F�cUqZ����_�B�r�py�E�Ey��]���Q��Q0Ե*H;�$l��"b�ϥԵ(
BG(��'��,�)�\��$���Q�WH���@�����f�.7�C������\�+�v�wdH����&�Mp�cLon'�̝�B3�=�j)�	�e���>��ۘ��Ybs �2��V�*� ��ǩ?R	S�����l���v�I9���QA &�c��5����S�C�f
6E2 ex%�G�x��]����r�_���dBSwj�-|]\Y����T%���d�S�+Eyn݃H�Y���K:��z�x�VMm��Dlt����|�ơ ��Z�QN�����8��?,��[~����iV�9M$Wi:}�Z�>�Rϓ�JK���ڕ�M�֛��{�(�{���!�l ����(N�<$��7�0�[j�)�T&�n�����bOd��h�^�&'�Ǹ0[(AIX�/0_������qy���bMF9�m��*�!�0s�w��\�λNP��"&ɨ��������:�E�aY�\��j;%�v�/\����E�d��%�0N����#+(�E0Q���K`�ݰ�<'wt(#/����0"�Tv�w�8`Sj����e��.ImR�jYzؗaD��f�(��)j�M9~�ԥVH�²֣�a�b��t�/f�l��8.;�E�6�����қ(��O�+z�o_����D��Ӊ��&�t��E:���n�1���ƺ���7l	��X�0�doJ�o��٦o��RVI��P�,����ڄ�^�4Bd�pu���Y^��n��̽25�i̪�!U�W+���_)��C��pc��r5nX�l���n����LX_�]�i�C���ű�=�H8	P�rY��'��ٟ��^��Yb�93@8+�,��I�P�I��X��)K�9��Nn���ZT�0��L�dg�o� ������v�����<�<��� ,��k!�,GCLADR�j"_��z��ozؼ�x�䥣�n�=���_��u[�p�p'���|�$D��z�Msg��dW׶tG���3{cm�ِC+Wz�ng�J$�P�	�)r��5�hR�����.��D�p�?����+����W�����~�u��&"bs=Â9�i�v��`4$=����:�z��8��n�$�~�+�ba���4C�j�WE�M��`�K��	s��鵘�3�t�����-7�Pз�Y��Z����U�A1�F8�W�R��N����z��9+h�Å��8����1�tI7�V��ok���'NV�G{)�?�mxFQ �L떝8�7�NU3��-j������`�+`�|��p�Z!�Fw$:�sQ�׸�!�-T�߂��ҫ��S;:�N�d;��t�$(1|u ���l�Ӵ�&�7D�)B�^�nx,v��؊���1��D/Q�*�g�6`�D��es���)�ш�(����F@��"���.$���Ȼ1O=d���$l�a�O���hN�i�{�.�Y$�oEvYk��s�����6�ls����½��-��<��Dt`�	��ɨ��p�H�at���NM��n���2�##��X�������O�;(�I�q��H��`�2[(8�P��'o&
�e,V�@�Ł��2t�Bs�P�	�\�<�+4V�f��֨%[�m����nRu��b��t6�{��Gk~���/���>���4���$b���zX��7��f3ǿ�i#�*vot���c���R�.-�x�:u�D3�R�>�3�����T,|�0��� O%"ȓ����e�`<='/�<鐤	�]T-Sr����aŕ��͐ٔ����r�Tks���WbM�j���m�rlr�)�Y��i���'�KתpSZ����'{/���¬ohgq��$��P�^#j�pH��K��Հ�V��,n�~��#�k�O�� ���4�{OOd�?g��ʬ�U��y��r�t� e!
)AE��
ƛm{�?l�M���=RhY����+�D]_q� ��������"�K̤.E��lO�wLF��҆n�*tj<\���S:����~�R�Xp�����ÿ�gL��GFo��ra��l�'���\��s�ΘRFSW�"��{�c3��<����?��M��V�z>�P�l�å8���G�Y1){�p���r,�A	݈�U�d߬�T�~�5�&�&Ó�Gu��뜱O"8���O�R��Ca�Y�<{�^��Յ-����k�"wS�����������#�n�ď�;���b�9��g$
S���(��Sl�~�
W���I�x�A#;�I�0����=��#�����6�/&��ɖb�����wGHK 8ט���~2������uRJ�b6�ͩ�&(a,P��8�l�+�%`=��,"o�
Q������\�%O�?_}���ފ7����_�����z���l�O�P~��f&��x\P2ޕ�L6M��w��8�A�:���0x��x�����Lk���~�%���3*���,�N,Gm��?��3�����I�n��)���E�6���]MɄ�u
�����̇V�F~��0;��T�0D�e`b�]kl#���e���˾�qp��ks)>�q�{X1������yf��Y�Jܙ@�O�I�PL=_b��7n�t���sh���<FC�/B���q���N�İa!oꁳԈ �RiVS�����-�k�{wS�����BAl<��v_ht��>�t�����8��VNmQ<mvMƜ��zOX-4c��Ku�w�+�N���}�::�wcI]G홭p���(��*n?ͨn����oz��E��?m�$ ol⠓c�~g�t�Ǵ�_#�{��w1�=x�@�M b=J����ɥ��Z9S�( m��?��ػ�oc���?T�y�r��,/�2?����D�e��G�)Z�8 �Ŋ�@�&h�Ĕ���|�tFR����W	���KȉC%O۱�������ǆ~�Ӂ��E�l�Useڇ�5�081N�kʮ'���'?�*��Qpb��_�fuub�Q#R%���9OVǩ�y�gHHIq���v"����$�4A^�)F�P{��B�?��K	wR��s}^�I�j������p|����v�1V�� �b��v��+�Y8�C��ROWޥ�y�[O$�5�5�k�Z$j�;�3���ʕ�2K>Q{Z�!��D�<�Q���4��%8�i0q^z�Es��r��R�d3�.���]�x���j~�i�B$��R��ᘈ���ʿ&��mi-�H# ͈"#��"=F3�F����Qҥ4�'ݍt�������zu�:?�7�#�����*�M���?T/����9�s�#v�Y�T�� ���A��vkr�,�2�W1O:��[���i�A�W!_��0f˒��R����{vcϽ���K$��)iy����j���(w\|I!�w��b�}7�'{Jv���$|W�ŉ4�rvPK0�y����������0H|�n[�֛���P=�N1�l�FX�7Ұ��vҍhl�ґ�T�� qg�B��%�_l�=�/���1u�ܖ5���2Сڃqf�VPa���O��-B����g��j���������7�$��m����C�W�}L�{������j�5�o.D9��N������I��l����[�9��Q��c�Y?`긟�i�{w���C����)�W�n�&�q����.p
.���;VM�VJ�bA"�*��%���[���쾲��vW���s����t�#�]�Ex9�ա]�	���r^��k�w<\��7���`���BE
���U�{>�n����/�*���D����?�����OvF�w��b�⣘|��ŧ@��(��GV�g��(Z�Ok]Gj
�1ՕZj��9<7���q������ �v��S����r"����#�Ι?e~�ڜ�"$����B�w�8HO_�W.�e�ў9X@��N����'�I&�4��B�Ǚ�O�]�X���6�h���+(�hm��ya��h�_�~���\0Km��u��ADp�y���/�_;���J4$qNr��2<�����h��)����H��B�'�.��;�brs��ζ@�N�2�z���`M�E�hL��d �(�p�d��E$�@z��"���������X�n��E�Ӟ��(R�Ց	�W�x�z���`Xȼ=�-��U.�� ����c���m�=	��Ǌ$�1�.p����ب1�"Iy��u�xo�������ҙÈ�1��tDB`w�T���a�u_Ư,��h��i~f�;�xǢ �l�r�L��Ƌ�3���T��V>=:��y����\��p��/�DnC��g�����y���r�����Ϯߑ��`N� ����p���kg�����M�v���΋�b��荎�'��R��~~ī4_E�)�~A����.�>�3R���l��t�o��/���g9���µ��H����t=�AE��~#�u�/`�:��v��D�\�C,NCW��~�֧*�ϒg�v]�}Db��茈���� 5�z_����;��|a������ۦG�1�1�m��/GJB�����`t�ح�[]������Ev��Ð��oMm �.�{k$�w�E@H�X��7_|��vۢ�IH7�{�E�ur��ڹ��N��iy�$7�	]����������Ӎ�!�����*���7;#�=22�tr�b��ތ���$>.t��Lj�:�"
n�ߞe�)��b��Ɨ��i�5��f��ڋ@�ʑ*s�}����~�z`��^$Ґ�G���s�TJ���-��7��iE�|�q�a�J��"Ph@k{��פ�G��]��9�g�TlL�UV6j�՝kr�Lы��C���T4�j�������!<�\�V�|ಗ�s{�;���LB�<���[�|x0����Z�Y�ص��yXz#d�(!��&�������)[�݉1~�wa�R4q��������s��G�H�_YjX˧wn`�9�Fʺ2�`Qa�v����U�������T�ofI�W�^1���	��N;��e=�u�
y���ͼ�Q����sx������xs�V����~�3�-6���v	�2��_,�'��S�Ȍ y�pw����ɠG�.W16��S��$6�W�:��FQF�>��Ynm�����*����n�F�b�~���������3��Dɗ�Q�ٚ.��+K���y�^΍���]佝X��$����dh}���4�=���%.��͙s�2�F��l���_
h�i�;�*p�<�˂�%�Ft�~aʇ�8�4E����hAQ�����9��G���}VS؜��E��8�v8�15�������	@�0����,4u���z��@7B?by��Nj<r���>��a� e�(xBB,�m���Y]�q��@�,#,�(�|�ÑSJ�]G�N	����t=�j6�S6�c ���fH�2�2FT�#Rهl�����b�W�
�����3�g
��GbW8�O��6>��?���ǧ�����r3�x�J�MHN^�����*&A��&���@�^�H�N@��`�6g�GhND_q����Et��9�\��[m��^�I�woח}�9ث'���� �u���cN�o�h�9����r�T� X�&j�5��~˟�7?/j�
�S[V��xL��J��,LD<o�@#�c8b��o�i!�_y§4f"�������Wx�'����"h~��gށ���ޙ�nH�`ycuE�� s�ٺQ�z����T�������C�"~U��,�'�_���>�{�d��r�1v���񏚩Utw���[�1��ߒx<!�ĥFZ��:�m�?��[�Cfu	ݫ�4V^hr�d�o{ұ])�W��wkf#��>H�ұ�9��J�fk���y�6F)c	����C��"�F�{����y�w�#6�$��>}��|�2&�����}�/�VÓ�#:��DK�|�.�	����װSӥq����՟ �`?�U<k�7�sҲ)t�6���	�_+��%��'0�F�d���q�J�_n6��,Sd.��k>�g�_s�_���r� �ל�lnY@�7E/���l��.:R��f�U�I�կ������Q_�9�hu��b-��A��n�\�l�Q����+�Ts��m��V~g�%����������%�#a�i./o������j�^+�D���'�{�f��$;dN�C��S�tL|�Ĥ;S\�N��)��W�g|��ޭk�&S-Q|SG�D�u�Z�9U&=�9�-(�fw��"��S���^V�?���_)!�'%�@/;x>o���x:>����"Q�F�q����ZC�Er��������R����J�a�7��V�?��N\�R0�1|�`�ئ�|��dv.��0��DS:�����5N;�B%��þ�c
��5�w����/�ӟ�c��3���E�繋V�8�2>��E�c��_
v�3��@҄�C6͎
9ڡ�o�7���:v
3S���a�z�(�Z����I��_R"1|5[WP�t���>��!p�ſ��H�Af������o%Kx�������������]:��h���ʂ���<������,]MΞ�C@�q	d]�-��T��Wɵ\#�!]����m$��1� S�	�ю?���
K��*�El��6��I���괇�q����đ����Y�D���_n$uŁO1���%����U�C�����uF�媬���E���jc�����^r��\_;S�Jh_�\j�7t��>�S0\{*�c�F��T���gl�9��N�rv���͒Es�_C�寤�X�����E����Q�_?+�ppd����P�!�6h��N���x�����$.�5'X�r>u4V��:�r��A�w �ȺǤ��gy=4�tʃ�	����91���m�9�&&�M�d�hp�CL�����T�ikcS�St�����m�X�C�L5qɨ��J�ʗ6�mv���ޗ,�<4)/hZ�ޠ@�I,�]�$ك���7@J��S~h���>���2{���d�na��}*����/[���0�J$k��:��&wgM$��LF����	�s��q
�!���e�I;k̭�H7��<g�1��)�O�W�����7M�J$�,��.�Jn_`�e��'M���B�J�;���p��;��Û�U�A���u⍹��퐙/-���_��}%��;~���8�����F���*�#'�æ_'�����D�^�a������TD���o��6 �I�NWB$�V����ƒ[ I�C��yc��.��_'3U��5�Uv4�m�g�m᥎Al�0D�~��hʠΟO�ѐ���n����/A��"9��r�#��.|C���阕,&-���⁐�%�s�J���B��&u�;��s���(��=�*�TU|ZA��@�ՐL�Փ������}�v��e�G�ؓ`�I�5��aw�3����liO��?ѷ3�M�Xӹ�!h}�1y��hx�~�e�x�X����.�	m� w�P��c���������Sy�S�:��Z��:���	��.���%@�!g\���09L|v��'~�2�ڨ/��<
S�m�*�M�D����h�`�_S�qs����8�3���m{ڸ\x"0��5��qϟT��o��|����=g�F��oH��<pq����&C7h�-��3�n����4Z�&g7�;��S�tÓ4)����B*�0bd�IvJ���,��̸���魑�w����!�~	/��1*4z[�\����I���.�����j��[]�W��]x�oZa�u���7�h�����I�~Nt-���ba�@�~��;J@c�g0�H
��B�����g>w���@�L蕟ч�=�Oo�^�#B���"�h�Y�)#fwRb��S_�Þ�b���G%�z�q��M�O�[�7:;�8 ���"8��<=k�q�>M덴���<��N��Y�M���l�߇HK�z������D�)+�PU�V-\yo����捯7��+�Wk���:>��	~�N&�V� QB���8��
��[[U��H%E��T�f�U��ME�
�x���O�(�J�y���7<�0<K�B�x}Q*�.�<��tۋ-i��q8d��pޝ�&��x�S�,��aZ����?�o�E�0�xoq}�A��D�:6uL����M���a�X�����ה��|z��]̛�P��!�o�"���v��X@b�xm?7Z��m�>�{EMQ�=�T���Ť5�j�C�&���$qoS!_4f[�����1���<���k0]�L�V^jʅpG>�r��,�%L�������1i�̟i�~���VSP�r�-y�؛՝.~a�/w��q�v�����0��1A�<7ope��?mY�?,~��I3�c"�lH����&�b���Y�_U�W�f�=I�Ҟ�O6,wH�:,��q\�;������c�3m��֛1�9�W�v4���X@���'�H,ZM�l��1���Ԩ=���{�z���.�}��pqS�oO��B�����vs��y'���Ys�i�7{�}$Rf�Db���j9�w���ܥ����I<)���s�A[�8vqR�3�\6�*^DR������/%e='R5#��W�}/v��%k2�Lmr���dc��k::�x���QU(�c{�Ʃ� ~�J2�?A6�,Ӂp,P���J��\��XH���۝�ru=�3zqq�UW�+����Y����g��.�j�I�$�O��U����+Zۀe���W ��O���]���lH�q���{�F�_��l��܏SoUPb)���N2w�����o�f���+���(Uad���Z�g��o�����i�]j����wOLC�������he_�!&ó�nҘ�{�Հ���gq��8$g����~����6h����Ԙ߇c\ u2+�%�ȸ��5颁�z�ݎ����������s��l��³+�pr�)򷸃��}Q��#{j8���~�����ɗ��LE\����"���C4H�YL�<twg{{ 5.ܖ�:�sm�`?J��^ѷF���	��V�iP@��|+�Bp��x�7$���Ι�v�W�+����
�<��9l]���x�h3I	ל_U�dx4of�ݕ��n/akÛY���H8�TcsC��O��������Uڣ�B���W9�F�#��.������ܶ�m
�mKF��jc�X-]Y���j���ҹ*� �{|7}m>s��,p�r��P	r�0x����Ҩt�:����|&-6�eR.wJW
�K^��v �XV���/�\9�R��Q�խ�J���U�+ye>#&e�S��&���	z��V�%��ڂ��6�D����"Eل4�����+#�CGZY����D��h,����Ё�����>U����.0eIz��:sjvV��
����rqQFW0�� h��; =��	wd�g}�>��='!6��-w�۬M�k�:"��R����jK(+-)�o�Ȳ��H}Oy,:���^*�YĖo��)�������M�nk�gp�Ѧ*�x�IJy�������n�%��������0�]��>h����w�wG���-}��ć~EC&׽�?���
�H�V~�Pp�KS~��3�N��찻�����y#���|8+��2�A3�
|��O��*��˂\?�T���J��;�ZZ�I�=�7�-�1\5)3v���fT˹A�'
>���V$#�$�{�<���l��-O�n A#C���
'4ȴLC�A�%y��V�+�|nm&`D�Y؊��b���P��E�ʬ)Nk���\V� ;-QA�\�Y�BL~"��`�/�L�-=tz2�{|�à-��9s��7�����p�<�;&�SU�]�h�e|9L���	�c*J�3�zqW��h��m9����P������Dͫ��Q`��A�Y=�b�].o�Q�Y��_�y�%kbK�_ˣ�ڰ҆�r}6�6��w��z �\<��PO}&Z�����\]v�5_�����ݼ�~[S�J9i���ʖ�C�2�M_�7��&||Cհ��u���k����Q�<a�T��Z�zU�$�
���G�h��h��Ǳƿ���nD��Q��;;/B*6t&\��9�z��:�uuT\�'2-�R4q�!i����k���w���}���)��`�%�K�X�Ѣz�X��6����ʂ�F�9ڋ����w"1򽾮���y���!6��{>�fY�g�n��#�ڮ�w�o��3�G��[^6����l*�ܱhJ�&��E�d���]m�G?0��(�δE:+<Zr�N�JEA"c���t��c��6M&L�oG�����$q�ȝ?��K��޳o��X��X�T����lK�����o'�T�t�r��ܚ����ʖ�D<�����<�ޜ�	��@�f��Gbx�]>�u4Δ��c��2�#(�1Wc�ߧt��VR`w�dգ$Go���&�%���IU�O��� �A�x�})o�W�a!B�Dl�����)Gcߔ��ň��S@�|i����m&�]��&s�A��R���Fb[RW�>�#��R_Z��Ju�9@F��j����|� �|��b��*.�ZE:������r5���8�<�Oٗ�QҪ�˸w3������QFM�H����d>HKF[)��2D9���6>ij ��r�+������e�x@������#bb/K4Q%��$����ŕ{��b~������p�ϐ�f�v-��;��mG^c�d�3ʚF���;�f�igv�&�-/>mb�\�q���-��[i�;ح`Vx'�_��ցE�⡡=��+J�0W���&���iqW�_���0�a��C�d�I����6�o��W�b�_��9�/�x�+�p�O2'�^)�ү�c}�d��3��n#�g�+Nne�L�qX~J�)�p���# �ߔ�X�M��)�V�ҩ;��M|�j�����/Λw����q�Z��-2ע�����$2#
�2EX��H~-� ��}�$g
I(Ȥ�-���	9��SZ�h����f�Zw�	V/��������#<1�j�?j��k�����LOS�+>�KF��b��ST�秤J/&W�=´DRNT�{���G\��p��8�%\�� �8�܎��1�QI��KpM�
l�6Ot�9��)����Ї�XЪ�~h������s;@dl����D��P��+qp�;�g��dA$�HͧuG_�1�ui�ȏ(���3f��\4���'�������]'���D|��r�u��s���]os#rd�<�]Z��eU���|O��4�,���[�y�R��r�����Tl����u���=f��V2�Fe_e�Jث��k�h�wBK͸��N�m���R�'A�hG��;9���*�r݊yF5��Ҽ�oȬ~��5��bV�B P������w��Ոл�cF/P=��(5�)��<��Jx��N�bXHq�j��$${���I���qڔ3���ic2�G�;]^�8�_I��[�eO���F�L��Uu�^QU���Q2մq�XT�L�-[j�����b=N9��/e�~�FI���(������l*����<�xg�g�Z̤t���9��3�w��ޠ�'�)����t@m�~(�?Ĭ�g������ư;�H���t��+���ty��v,�Щ2��<��g����sL�J��w.�`~-[p����UF�(����j{��y
�qX<�6�ǉ��?r� 8�H�� �s?
^J]����� �Ͱ��C!�Dƣ$SAV�c����M-<j�T���h��y{�8Tx��U��X�󌻿�O�,x�k0&��W���ώ�q6Z��^��Ή�����p�����6e�����z��H����������N.�Y{W�_rj{z�ΐu���Y�m�2���|��S�U��۝S��}��i`u[�������֯7�)Z~���S�I��?�P��c6K��W���޲ZR�f�r���2����"�2�}���,���K������Ɉ�E�ꔩm�b����׷)U�ܞz5�F2_����I�7Cʄ���`1�{c����l���Գ]��lR�E��iۥh����s�_��PO�ZF�.��\��O����Z���6�5�����\M�}MN�.�����H���u��.����F�_�;Swoy���_�c�ѿ34��5�TdKT���K� ��N���_�,������);���~�/�%������ ��������Ų��B�-�z���tks-����BE�R��PK   5^�X:u�� �� /   images/3d480ee1-e9cf-4ef6-9de8-5a7043d7f31b.pngL�UT]n������6���K��4��ڸ;AH����4`��>{_�1�j�����Q�t���1(0���UU�zpp�[pph(�WR�x>�/��z� ��Y�88:8U�����C��������ޯ���F�.���z|�TM�Xϔ[����$?u��@`%�7�Z.�c+<b,��x�I:�U~vB�������JAN~�3	y�f��l�g[�3���-	�'��䢻=��?/�fߊ��Ǵ�2�2^��/[��QG�jj���k���������Ȋ�r�ۅ���_���;�r�qY�d�>{4U��`��	w�eI +���|?�+��6�)AH�D����1l��]Q6��8���y�&R��zF'D�h̍��(;�a�/�����������}�6�'((�WX���GcM�����9έ#	P�I����"�=\�U��LRct���[��?���IE98L�)L���C�����#&��ȃ�qY���$��A@�K����'c#i����3��4S�Xa6�ECGAʯVP�#��H϶��n�`�,<}�5��ϖX��?���\�� eZ1\$f2�4Y�Fa���;�0g�y�X/��\�J���~m����.]"�<����1�)�k�l�Ѡ���_�-=@�!~�65�s�����q�.�Tڜz6�,-΃��L|\�4qE�$bV� ;�`p7���c�A�ƒ�N�-�����>>2���C8�>���2�O�h.��@��I�����NG�z�;*LVI�����(3ނ��me�����(�n���g�+���ռ��m��ni�n&+����N�5�;���~�.��$=��6�=��f�I�J�C��/S�}riD��S�	?C'��,>Z$@����Y���m�J�A2����-"�?�]1jZz���1lE[����{���=�8AX(�
���	;��^�|X}}�d������,��G�mf<7b�~y�;�Ɔw������8�4�Q���s�/M3-�O��\V�$���Po&0ۃ�D�� ��Ҁ�I�Onf(�_�Onw��0�s�� N�|�Ի�S���C���J���a�Η��`�OAP��ce{���䭞=�E��4�$���	l>�ehX[k9���@ݲ�X�',ȅ_���<�U���ٝ	����.�H �H�(���l^����+��`Ҍp�����-��G9Z���|�5	�܊UZ�C6�V�@|ُX��@3I�L��%��qes��^O�?0�K>��� �X�Ak��lh*h� 1v]��P,$~>��;ɮy/����h2l�y"�T��.���&�Cң�#/,
|[*��B����Ԁ� !
�ua�Tx� c2�y�
:�'�]�s��⏔��2:5���CVz�,|��ß�+���G
��~�����˅9븄��������v�A�H(ջL�
\�t���I��^�=4�}���x	��o�F�l��>�?���~�P�Ϗ��2�Nv�U#4Z�����<���5c���s�9t�m�{��X��b��.��]��0,����2
#E���,x��CI��MTHY�,��`{�������#���b����}ި��9��?�Pf>�I���
��������F�V�b��~��k�]���6��H�<O�g|�.�2���@A8&�ȉt9�kxRS9��_1��x���>�69K�{���K�����^:��3R푀I7�cD�<���Y�F�	�wk�����!��FY��� (��o9� 1�V�'��P��ڇ�>��p��O*n�ʞ�ik�a81��6*
(?�8�iV'5�<.��)Ha�hMRXxF��U�g|�7W��kt��"��J��_]�C�c�D�t�e?l� m>e<�_kT�3d	.���u��s"f*]��1��-�:ur��u
��4���A9��X��+��+�d�ڸ~,<S��xa䖃��IN���N"2��:��~�4����w� �������o�/T��V;�-�T<����xV��+�G�n應��D<[�|�[s&�H���"����r��A%�;����X�H���2g�
*.��N�YlY<r)�-;9>c���V���-3&q'`A��̉-�/��|��%��k�/$"�u�����}�j������e<��}O��q�kO��3�gVD��?V)p���i1ė����=�D�2�!�?
��U}A�D��:�g}������@�nz�|rT�"�B� ��X|Nj.ǂ���3lo�cQO�E�����BPP6=�&ⵔ�����?yT����N1��B4�^�Jo�������b1�%R���L���^��}����*kޖ6����a�?!լx�Ji		�4#t0�X_����������F�����L��R�n{�ۡ�����7�P1@��"^��6l�ŗ�#.��0u��8T�4�0K���u�I�?�#*$6��t��[���d��;��(�A�Ӗ:A�"i.E7���TVV��!G��5��y�q(�Uq�`�Y�l��6��\�%�L��eS
�'����m.���գ� |�e��\.�,�����?�(��K�Q�+]r��W*�?H��Ǭ;
P�A̡�	�Ob��&��x�	�'�b~U��`1Mj�=~<�kҕ�b>���ؗ����9�Ė�N�Ô2���>�����.'�K�
m��7�`(}h�j�f;�	o��HޓjPd6F��B�%(l�FS̔��8n�[Rc�d���p*�0t�"_"9I�����и��p�lZ�eǜ"-�+�*�p���
�3.D�#�x�/���Z�4�PNէ5�a.�q9����H��.�5\��:_�B���)��y��H7��Q�q�8$��L�e����ĶդSDr!��>$��ɁW��菢���`F��z�%S-P��XA�(�f36��� ]%�<V"�����K�dr����.H�L`�y~ńV�܌���b�C��j����c��agOo���d,���/�w�^Oh��	ko�z���)�8A&�N���ULR����:e,��7��F�M�[9���ƚ\�~�@�-���Ë��d=��s��(¨�F� Zga����e��0��Rs��ZA&�g��M���CcZ�:$��FR�(;":�G���N�n��˚���OH��Ks���;�2�E�X�Ĥ(�?58SdI ��/���t�
�(�'�]ܥ�pq���u�Z�G)�����"���w�4q�j�.�����!��i-܈�rcCi�T�g����L?-K&@}O�B������T�j���6%���QH*bdE��ɆC#h���a[���F
��҇$QS�P��a@���m�^«�ӬD��ԦM$�*��'���ŇP��A�xq*�h���T�R' ϐ�+5��#9=�N�1^6a�yv&���q���$ۢ@�:a�|�eH�D�%��3?���7��؂��G*�0KL��fL�B�р����?���F���G
4�=+%�Sp0#Ȝ!�!�7(T5ub���n:f�D�����@Y����ۜ���L��ot<q��A��� �G=�����Ac�8�r�ّ`=�ŗ!>d^n4|^��[�k�Yp����{�`վYj+GH!e_{y	�,�����%="��	y��T�%�i-	�f2���<�]�����#nSL܅�.m��X��7U��/�����a��b�TD`*��Y�{�b����H����7e�����2���,ar6�y��d�JC�a)gh�
yRw��+���d���P*�A(��P�
��T �8�!�*�	�-Ω���j��*��&$y�  y�!�@���D$�:�i� !����8t�E�T7N�d�MG�0%*���!�$���m�L�7[B���hl��1����6'�P��ĥ �f����65K$���&�H�t�PF��Ț�#t��n��8~<��A^0�r(����!�zzl6�^)�}F?h��r��D��o,.�)fɡ��Y7�^��6�i6�RUb���V--�(1�0��+�f�J�!��N��y�^([BZ����Fa��ɩ�t�<G t�*�yi,
/��b�aHǰ�n����U`�~4�CQoK��πo��g���V��`Ĥ6wFK�t�����h�����TS���[����X���J����M��z3�O�\cA4$�ػ.e�OZ
�����!�g9�oR�����pk�-.l7s4�W[z�Cw� a��h���)�RU��&�+FhL�6�b��G�D���/��H!E���O�qU����ٖ��t .:�v�g���L�j��x�c�db���5�?�����\����[EJ�xmل�I�8�"�p��T띈Z\�>�S��Y^�C��B~<޶]�0pc�)�R��WW�$�����R�V|d�R\����S�����ሺX�[[!�5��b�?�/�D�0���'W�)R:L	!��]@�H�tG+[5�
��q1�5.�����[]R�&(wB�
� Wn!W�a����Ĥ7|�5ΫI��l������A9D���l����q��/�"t��*�c1��B1��k{?��ڥ����H�_�����T���/�Y}Th/���ό���t�+'5�c�u�Kґ	�;��{�-�E��Jl�m����SE��y�a����؍����Y`ݠ�_S�J��`�!�9� {E98ܻ.�\^^��k��Ff�&���R���j���9^�G3�_k�@�B�H��ܿgt�������w
Eb���k��T�1���Dc聉�6m�;�t�2д�8�r�z�����d�H+�Ac��~`�6!�s��:��$V��|ԯ˟�����gw�$��S'|��~��:z�b
q�~4�H�	�ZyFne��6���t��>�3?����7��CW��xj��At�;��-��ů�l�T]*T��b��'�D�}8FZ�\)�e�M���p!o=���=^&|)�#N�U�LMRR��� f�!��j)�^Y��\EC�D)̎%����A�ė����ē��wC^��[�K����].�y?т�,񐬻�CGO,��z�/9e"�n{��$�y_��:1�A�D�U�8�{|EW��?O^ ��ď���M�K�e8h��͋��T_�l�Iks�~��*O����|xld��)�g��8�%�@��ֈ�icDU��F�{�Qri��sH�i�	,�+_e�Xe���r�KWԑ�A�#�`F��%X���D^D-겪��Om%v�?�X,�0u1�Jhy<�7����@�~חJ���
7��n��Dn����}��7��� ���͔DYV��O��1n�$9���5����bH|S�Tߘ?8!�-)�SJ�T�4a��Ǉ�?�hc2J��c���"�=�mO�0��b�J}P,"9��-=�х��ˏ`ч�1F��mPZ���
o)"��~Pc���KX�j�?�����mfsX�mqM�u�X��f�c��ʌ�N��(!�gԃ��T���1׮\��c�@JE~4�	�m"Y0�E$N�o	a��)���aw,K\�&���-�W_ٿ!*�@Y+��I��m%��⿧�5'����Ⴑr�
�~�x�a��l@<&m��AL"*�U@�j���֒쒙`5��:,��1���w�c�%�>��An-�S�#����IMjH?~ĺ��I�%��]��d��U���b�����,;}o���Bv�o��mR�����_��N�ΪK9Η�*y��"�2N;"C~B"�dN�qC��Cp���9��:�*1�1��� ��vuq'EF��~�/�@������=r~��;�����Q�4�� ��&CC��2�0��T�X�/R�f�I�����J/�&�Vͩ�Vv���t߹js0,tdG#�����mk�p��q�C��a^]�WK�|����"�n�JMRA���D����O�ĉ��܀���ET%�+I���@�6C�k��`�S`�Z�2jۆ��Ce��>�R�DA#]�?D�7{3�ͽ̤@Q������P���4]�YO=Z>*b������D�����k��X�P�sL�&i� h��X�͎�_Lb�"�Q�:�2��O��e�x	j&.��(�6�$W�/:x�xJ�_=<�#-E��O�&��ۙ2����k��O$��B����ǩ��M�z���Z�Y=z�� )���8�$�b7NY*�~V�UL�Q��O�ⶨR.� oUeuMG�O.j�[-b��qX<1�h�O|v�v4�·"+�e���{�I�*��S�s��֞��48��ȮL^�!�\�+ӄ~�-2q|� ל� %�\�M�Ŋ��Be�mce���d_3�ÕރD�M:3�!�4�iTR� �ӈڙ�jeD�QZ�<{�2pf��g�~�yȪuv�1��s��\?���si��=���>n� ��~��dE<&�*o�)�
�'.����7{��Y��y4=O�cٕ�=�C��.Ν�(�
�%-��i�Aсˎ��ʈ�kA�љ�»�wNß���=�@��1t����Fz�m�lQ�4�-�F�H��Z2�઱��*�T���c�$+M�l�>�h��H4�b�l.�x�tﶷ��}�:�"`���5��JP��4������6+��3�?�y��ىԠ���aF��(*�u��;=8�US>h(I�-}Ý�r�1P�0։�[�M�h�.�= �↼�V�Y ��y9,u ڡvZ�^Ȧ��d8\_d7{/G�.�'ד��`�à (�6�V�R��(����(�����ȶ�:�Nȡ�GBp��&7 �n�ꌢG��'��\PS%�WG0Ð>�QA 2�ԣ��C�#�#4g����#��$�v:{`t���,k�OD0O(u��Q�b�����j�FV��6���D\v���6N�7�<�A�a3�������QN�K:������H�����p�H��7U+���O���
	�^�����@xT�H-�����z^�
$��ԋ�S�9�,���K����F	��
�G] M���'��$c-���md��iP�4҃��y�/�����(X���Kd
�t���PS�ͽ���'�~����)��������:�C�dq�x�<�j����CY|�P��-�@�fu�u����C.6d[�w5������EN]� �F�&1��3�N����L͟&����B]�CXw0�����>07�x��7�Y�gL�Z��|󵝚��j=�nJ)ZU�@ٔ㷔~�Ď ����#���&��=x&�،��@g�r��'IQ��п���߅4Q��v�=؋�f��Cp,
�NF5g ����M������B<bt�=�W���0�f���2b�!��� ���������u��K�l�#����3&��5�-Z�����5���&;�bnV/�_��#�[�PS�U�Ym���	s�(�o � "H�)���������f%��� t��}yҐ���L����Gm�D�!9j#��Ԋ��ٻՖ6�Ĕ�6hB��`��S)�=ޢNk��do4�a��%�)Ę����������:���\�Ng������X	@��q�����
�t��}�zR�o��%�Ѫ>�ۍ��C�H�9nʐ���h��a-7s�<dKA�Y*��ֵk�p�p7P���x47����.����-�)���q��]�?pv�eV��ҕ�����%*����zN�l6dފ�?���e#gs$�y1�*��)�|C9�;�{�e'�i������S��:!�[Q����i�
�{�<�-�&a�[���͑�N.;�T3^g�n�l��jM��,v��֩N�n�t���׶�=�uoʌ�S�� %�^�8��d��CA�QX#Uru㢕��w3�T���p��r�0v##�F7�6y�&t".�If|�Uo�!�t���1��+Q�H����U��f��� nh#L�� ��x�z'��X��{�)�g����;�T\�y��c��Z�'��L=�Sŷ蜜�zD��;���1��7jE��UK�����V/�g[��!�����C�6��1���L�"u��k�'W��9 	YM+(���\i �͝�`Ū�` ��>��u���x�^��rP����.�e:�XL~��eF�G�0�0��Ѵ���F����Ʋd��`!%$M� cN	~Q6��4���I�!�~H�,�X�D�M�x
Һ���5�� $R|HG�@�+bӢ�)F��!�pfVz+�5��U�:�> F�uY��V�:E��0���Ro��{0W(��'�(f���*�x� h�=t:ǂ8�r"��2ژU_�8.إh�����!�w��zF�%C&�i�PK#�V��[�uY��O}��3�Ă��S��h�t���&+�`)��Du�_�){�����(��3uL<m���'J�Yy��x!����ō@{�S�e��)_�V��Q�p�Fn9B�x�PQ{���չ?�wasø����,Ԛ��G�N�ֺ�]��U�`zB��|����u�&���s���p��~�s�ң�ϛb�Դ����3%�ݭZAA"6����IM"j��K����j�e=�v('GÔ(��p�R�xG�NrP|�jI�pȯ#qoB@��ӶB�+�:�b�A<
/�~��q;�i�Λ8�~-K�82�tNԣ�#��FG�ӭ7��|o4��rO�h�}:#a��5��ih7e���fMu�r��l��X���F2����[d��<���%L���{Tl�F��M��9W����z�ſ~��r��4nK���
��nl�?��>,t��[����������ܫ�����2�|�'��sAآ�l�!�<A�,v� A�;$~an��ߎ/z�lNP��X-��lL)Hz��ПsN`/G�o��G!W��Vg,�.g#�줢�������]ȵ���8}t�{����#��l(�竮��wq�H|�5V����Qo����0e"V=�Lzf���]���P}��X��lܺ���LF9�ݡ��������V������
�D��f�%9��c
/��g�Oi�Ոﺜ׹I�b;z����-�<�d5�g\�ҶL�%L{1��Jq�
�P�OrF�NB#Ŏrhci֨�L����:��&W���W�0�c�h���*/�C1�R�&��U�%/E��>�K�%9�7
�xu�'�87 ��1�*�F��k�pԇ�C]�Ouy��0���7�oaO��N�J�r��"d��7h��
�gI%hDy��	P��`!^77������YH��
y�M-k���� �LW��4}�!��� b˗�m��^��sY�߿2��Cu��	�j�\�U�$�|�PA�k���R%�!�{/�D�tc�/[���SА��WQA+z#�t�qX�|��~�\7]���'�Gfe���xA�ZԚ�p'.�m�㇝Y2��J�#t4�5���W�6V���]"*��
�4�}u;�XR�yuf;��p9X�>i�������x��)K��EC]�ʍ�G��dXuO��5�W4�J/�4�z�ɢ�x���b9���7�<�R���1�\�]�N���&���!m�C��jyv��[� %}��&)g=?����I�>���&�#�Q���=��fF�!O��07��K�Z�8�h�YiS��#cq�/�4
���Z!w'�%����J���	yzfi�⸡а��Ȝ�5�D� ҇�>1j�2vaX���8.�L�,���EP��P���Ń��Q�n|���N�a5�G<A�G�D���N|3�b�皆��0�J��?�?�,�ZH%�b�\��� �~t*2��b��:Λ�zkoC"mo}L暹�o�>�7�tN��6`g7X��e�ח��9� Z&w�;m����ʄ$��z=pn��*�\����F��5��C
�̚��I�v�Ě�-���'yE�=������߼�f��������J�pQz�)�d���z�e*����P>�E?�Ky��֥�`��y)��58�Ӂ��dW#/�?��ܯw�a���Ia���+�A�#����=�ϙ�̮3����%&h/p�n�nw��'Q.���4H��J�BR�wF�7:C�D�l���#��	��/+�Y��r��(̴�#�4	�jD[g��9X�1�Py��B#*��;C�Xnmȟ%�7���I}uwMZYCJ���qCZ�JV�v��:�Tx�.���B�z��(�,t2C����F���7�\�J�]�l{Bś޽m19��EhBMG�U�T?V���y�����^2v���YQ�����`�D��[fV_�	��S�A������' e�˫8"/e]�y~N��o�L�8�k�!G>⤟\�>�8�XeYBG�zԚL�
�% 9����L0f�4�[s��[ӠI��U�s�D![E�O�F���co���s��tTX��}b�-�P��jv�ڤ�"�p"�+�#���aY4��w�(6~KN^rrHF�&a�j9�/Z��k�T6BT��j�Pt�����lR5��ޓZW!�=����O@j�K7��f}���"zD���/v�2� �+2}���8
Q)_l�fitd'Q�P"j��h��g\ʚn.���ڑ����U����8lcg��/��Ha�:dy*�Ϛ��boa���A�Z5 �;Y���?^�\{�*��ęvr�3%��Y��̧�w��yֺ�;��B�ލ���F��]�@���c�
M�j GѠ�7��̆��A��!u�b�-&�LWa[>����$�վ�0����ۥ�MիF�o�����έ�M�?c����;*D�]�>��n!�n��tlQ����7k�H|oWwu�%%�(h�C$y+�ܔ�%r΀�pe\�����ļU�r���0��@gm�.��J��b�m>� ��B�V�jѹ�eG[���M�IuSD=�b�\*�*�D�tWZ�cM�U�~�W�X���t�.t�����*y�@�sYt>2Ъ��@[��Gk8�_l7�����ˁnq��!��1�D�U q�u,�|�c�8�ZWFv��o�3����ȼ+%�7�LZ� }���.
��:�0�P=ym?4F���w�nc�eH-����A��1&���Vc��hE[^��x���t��ݜ��7�V�?3�7������KO��p�Ml����8�+ҥȿ�u��p{v�x'�b
�9�=Hl[1��	)m�;�c�I��F�]Px�g�?۫~�����	�0�������9`����`PB�α|n>��%$�`��D�:�b�_�GXe�{V�W8-*�T7S��isk�r�=�X�n�6+n�x���8�'������A�W%��Kߏ`���`}�G�|RtH�o�Ԑ��]�^G|a�3`٣ ����~;/}���;���R�H����� ��8@��.r]���g[�+��x��2R�-S��_�=��C�T
��F�����"�D12�8��ᕾ��:^MV�"�ce$S6�i��(J�};�e�^��bx�^���dgp3t����ޖHEHa�nC
�i��Ku��R��*$;�3ε��_M��t����bw�e��Q<wƃ�o!E�,?��î�?�$��|��f �S����Ǎa3o��x{��bc�&y�1�6�+Q�r:�DǽzZN�����;�L���Y�d)	�y�������bɟ��kuć 0�隺��<������G!��U*��὞�rF�� �f:���;�����i7$|4��Nɶ L��}�2��G#M�3��b������)�"'��EM��C�TW/�$��Hk�a�d�g58�2��>^����-�xz6�l �7����oq];�N�<ڻ�F��E�A(a�	��+�}�v�������ET*��C"'�h$F�7[�
/4;��4���Ѽ�jBb#6H�M*6�ޝ�hl(-�$���G<��@m�qGc�����3��s�x�8(/4Q�bG��#�>p��3E�ۊj�d�)�
p��-2�b�}gg��@�E�����!͎?"�4Z�Ua}qj��(�U��i%N^
tڈM����>ou���?YYKQ	���[�-X�m���\EH�@�ҽ�Ԩg���ҤI꤫銥1�6��zǥzt>��ªG�$�B�'�΍ϾKFҝC"�K���{	��J{���ѻv��H��|
�+г�К.׭�0d�LG#����y$C�(�%�ǖ,��^���Km��ۚ�Ŕ\����q��� �Z�M�TYFj��C�O_'����q� �sf$S)�;m� �sZ��ө�T�m�VO�^����Yșdu��r���t�����3H��(����h/P���ۚ�l�z
�lc��l�M���W��z8?��~5�u�a���)⫵�u5�C_��4��M,�:�F�j3@'8i�7�5����Ǆ��-z���.��V4E�gV?-���{8�m���C��2�A�Ճ/��T88�d�q8X)4 (��i�P��hQ5:�^v�/��c���52�{��f��.�c��_r��u�Y��j큉,�\"��C<�2S����)��WI�A�6kW�T�O�$aQ�+gT��j����v�	{�18 ���ҽE�M�FCD�s>}������i)�������:��)������A\gY*[s�����kO�?j�^~Ճ�:���V��6V	i<����>�	Oż1������@�Aӫn�O�)Z!�SZ�V����zO�f��T׺6ֵ'U������7_XK�1X�ǎߪ�I����9|�R�K��Q�a�1"���6�V�	��X�����7��}��<M��zS�Q`Mr����u	׵��� ,�+�_=�A�h�U$A�0D{~O��x�t��#�v�ջ����3�����ӇO0�mhB/�A�0�zG"�/L+������h3y`�ˢ����OD�k�
�]�r/hZ��rB����>u�:���J("���ELZz�C'A�-�^_f�
F��a�o-ڿ�OYG.�O�[�X[^̸��d"��ȩ�kWWlNRp�jI���E����19�,U���8@�8c�����>_�B�6L���s(�
Cѫ�\lmC(S�(����m�?����ʷi�l[鍐���}�1��,G����+'���%��3�E8��m�C�Q�zo:<�wpF>�-]��@�78���@�
�1F+;|��~0�Y��
7�����8�3e�H#�Z
��ǾS�D���{���
����vͬ���j��� �33F��βQ����s��/�s�9����¨��e#�mg4������*��VA�*�p�/D��`T��E��Eb�|%�C)�Eęv�r-�_e�V{��5�6o������'Ad�P��"oH�M�Y/��M��
u��O�7B���������o�A�Մ��z�n����;�a3Y�^]/�,��������.�D�C�����җ�� 
��4}X��$�{}��z��;fo��;��);kW�� �BQջ?uj�ZG0�s!2����j�L���	���z	�r
�������3�!�2�-�m��/�,҂ɡ<�v�N�t�"S5�K��T�@�a�K��n�C�!s�#���b�A�=N&;��&�?r)kRč��	��:^�so�������v�h���r�V��.F�~�������an2V#�'/�0�k��:����Ɗ5����)��ko����W���l��N(�]�N��Pf8�ɩ;�=_R�珠�5i��ȃL����w6��l_=�bw�=���6Z~���㖛D��*��fO131
)���S��à��}w�i=�=ӑ��K��xc���Kӳ&Y��t�P��{�� j�gVp�f5�����M1֠	�}�6�+�Un2��J���q4x.B���:���j�5D�\�aY<Q���!ט�(&J�)���s�%���:m����`4ͪݕD����9r6g�,84���D�
��������Pv�@�A~ݘ��2�Js0�����:���U�9Zm,Si\�I�g�����&�ђh�`����}N��JԂT#�����>���M3�|{&Ã{�t��cA�K9,"
j�y�i��a���l9~8��#�7�G�s�c�uo�u�k����{�ϘO7
SIX[W�������I�X]<�g!2�0�4��*P�Y� r�ʽ�r/�g_��O<���d_ڈ7�~�`ϋ���u��§G��;���)������{�~��dj�]�m���i�pzgC}W�4������Ŷ�+��M��4@�X�b�BU��R�9����[l<�[���{�j���1A���8|^
1=O�n���Н�7��G���� �$�{��_�j�3�t
�H��kq�[�ԉ���r@�'$�t�F�d�����\�v�O�>�q���C ՅE$�,�A��~	,
/e����7[��Q�>�C� �;1'�&�[51+��F����3iؕS�z)*�5���q���Dv5F�0�\�q:N�Y�/�uV##���e��{��_=�;�l,���"�;B��i+�J#d~{���5�5��@��i�3	�9��ԅ�=$/
߫ �K8-X8n�%e��n}���*t��"0�14���L����l{������-�G����TK$�jO��.�G̪7eX¿ix|�	A�*���F[*�P��o�F���hm�a�k�3�������gAQx~?}�x9z�_���2�O˲��h*��)7?A7i��V���ٍ0@�T��k�\��&�:�"�]�'�b�[[�9.�M�u����]�e�=��pO bߞ
�rW��;�D�\Ҁ:&��P;���N���S�J�
�:ٺ�΍lܧgN,�Pfci��"He�DR.�J���[�DcS_;�)䵀=V��&���/TD���2E����?I���t$LU����{���P�jonj�	����J����%y�
���K����H:p���\9<�[�#�'��)3���оЋ�c��3��nj��%���{kI��B�M�;�v��υ�\���88e�G�F
�x�H�����g��z�q���]�����&�ew�β�D��!��-_׿�����G	��4UE�5�Hy-�
��'��̄����B~iNY������'����u��U2���mJy���N|��ҭܐ�Q��Y�tY����ÊQ��ac�6�0UY�M5��;�4H��N��u�e�|o��J9�(��`Kh��[4g����Q���
��S>�O(����C�=ʸ#G�T�A��&�.�{��WxtH6i�'�^�r��^�t��e�9H��F�e|آ:C\gp�	-�A?^⺷�n�D?Jٴ�#�_8��?�5o;~���-�'���*�_OY����?�6:B��U�U���P�8T�(�022�Il�ٷ�j�j��������x�@~)!4�Й��������^P�p�Z\}��ɝ�8/}Q�n���_oQ$'i�}Z����E˱����)�\R�G�p�ԣ3|t�߇9|�s���38���ٔ�Ra�aW���)`�l��nӃ)�{��E�������D(��(a��lLa��!F�G�?���F�KXaz���9Mg:v�|�o� �V,�����-�^]a���[.��wc��eؿ���A�ǖm�Ă9R8"����y�B:��\�S=�&cc�8�NT�y��S,F���xD�����8A��Y���ّ?�	�'<ﺀ�a���4�;��FE~�8�F��j���wmM�+����#��a����Q�����z����)�fxTs���YA_a�h�i_9A�v!^��N�!
��(�Q����^}.��W�h�sT��w�α5�Xi1r��LE�gŦ��k��a��^a�U�lя�Q������4N��6h�/�8@��/N��ч�q���~��8�"%ovz�=�Eu�O��|�vn��:mJ
�9
�\Y��n\����=*����h� ?V��Ir[x�7��@]����sC''���֔��wgNA'���m:7��ȷz�o?\�	��e�'��,��pM�8�i8։_�k�;9�ɻ��P�0����P�7��>�ɵ� K���`^����^1���g���k����/�$5��H�kq��ji�:�kȭ�������<�����w��Wt��9կ~W��W]d�b�s�Pg݃�uqp"Ny����^�@S9��U�&�,��O<��o��&([x,f��^�ح�R9��R@����<#��5�D�y�g��z�"D�v�J�\��@���yZGN��)x��	F�!��x�N�esw�"3��/m A�Ҙ��f�T"Hp�/� �I� �Q��8S�fqq�o�J��%N���K��xj?��?�/�v��CM�1[��,�X{���!
Z	5��v�aF�a�c|x����M
.�X���	�Zn��ʝ��",� ����!�6�w�4���@z�o���6H�qk�a���A/�:t�\��1b����&._�����.�_l�ݬs#��޹	9/�T/aay�k<i;>�t tcR�ܹx�u3�d��<���G�dʛ��S<��(����&���e�w��9�~�Ӆa�0w6Q3r(�氹��8�A.h��+0����Db���2�I������v?���8�X�F�-\��7p��7����4�Fm!3�{�T�I�3�67v����=x��
�a=��ZF�/ϡ��>/}&ޏWN_�Ƌ�xi��3�r�龰?��7:`NF���)�;oZnr$BLRR�%0PS�	�yL ��Il�NB;��i���6�WA���fA�r"�mt�e\��q��_�����+mkǡf�t��s����x��Ӵ�a"|����/EJV?
�|_V���T
G�zh���@
OWȠ�Ê�V0)ħ�㩹*S�_ ��#�����)�W�^@7�^�f��o`f���W 
�5`��H�K[y��T��MCʹOp��3H�R�*:����ҥU�n"��^�S�K.
�x�os��Cॺp��I���%�|�M*w�8J��������%N���K��xj�;���N�[y���BÓ}t��Y�(@�L��E��<9���L���S ���[W )���eD�Yn~��u�cx�=$��!�a�v:v�W�_�/~��p�W�i�m�/�ܜQ��SH�"��*�g�Y �j(l[��x�������4�UL,��6dCbטop�}�R����P��s�H���z�5D?���v�R��'��2�<�5��g���	�	��*���G�7�*P���
����
��zk��X�Ǫ�"��2�媷ZH�58�̥-���z���軐�	�N�Ϟ۰�����m\Z�Y�+��K=~\�9��O6����#�C�%&1*��-��\_E�Z�ń�*l�"0a:�ѤF�goV�MU1��yśA�fX�O��!HnQ/���/;�-���א�\��#?n䦊�^;�R5R���N�ť*���I�}�s�C�c�F��^����;�&��.j���]	�9G�����}�����,�LZj1����{���3=�9�r��ᆾ�7M`�@.�p���(�e+�!�a��Æ �0���-��a6,�a�VZI^H�ĴKr�!'s�ܹ�o�PՕO�s��}���t�rwd� $g���
�N�����y�waN�U��xGl�1�f������2>,�֦�-�*K����JfГ����#���FcfJ��Z���Wj�T��A����ݜt!����^�Ǆ�`���- �Z��Aο/b�q�?�>���`i�
\� mf��:����Q/�.+%*��� /�)I`�a!��ҥ53���C�vɵ/���x~oo_���T]���M��A*�E�2�e����b̜���x�����o����b}����m��xE������(;��F9���*���A��X��w*�ɕq��@���������>FH�^�
7a�Qc�i��VP}�	`��p�� |	������c�x�?�\�g��j���GJ��f�m:1�mJ��֘�\Fg2Ҍ�]��͛��j���_���!�gfq|r<ޥ�K�?7/7g���5^��+eS��ࢆb�B2�����!���~�e�\�����`ay�Gm�"
1���De�W��}�έ���.�N��T	Œ�:ӹ�8��ڜ����^��w�:�� �I?��7�����_����e�����f�$	ݾ��;o��+Ͻ(/��h>Y�_����.]_Gm�.��򔦬���x��<==�b�0�X�'v��8�*5�z��S)@�V�.�!�QqNpoD���	Ey^���kG��w1�)�f?}��w�����̠?��s���D���
T\fPz
xun'��+�vZ�q�K�uG)��g��*�x9�ɲ�-�Z ����b[��-=ֳ��WF���"Y�aL5��펁�DB���f�^��_���Q*�%����H軃$xͣ� �ߖo?�`�5���V/�<���w+����O�U���S��d�k/9u�	�{�R���ǥe���R�B*�K��{{��e�J�I2��h�z�|��k� M��W_}�?��������9��~�f4�&�f�Gf��x�����͛7�����ֹ��L���Qvp�s_!�ݼ[Ǵ_�F���P�wp����(�ۘµ�]���1��,0w�Ge����%D��Qr�`�{�E�u?�\�I<�����9��F��)��p�Mq�T�(�h7;(��f�P`�Eؼ}[t}����0�xw���ħ�Wt�zi+3�U��5���p�Ow0��ٕ��2M�و��DY�o��;o��b�A�wg0���V�9�{��\�Ts�q1;��M�d�B��\>�[ȡ����������������'߆㟠�x�F��1\��%��3��cQ��g�� �LעL�A����m�{��D�a'����z�ޝ[���\��]D}fJ� d#^���ycd����+cW�����=����p�l��v"�T�E#!�	I&��q��Ocj2��p��-4���}˃�5R�������[@�&����x��G)޽_�0�������>�e^���/��;}a5�<!�ײ��N���xE6�D�����خ�|�����l�]��5���M5x��c^��:KY�e�)�3�%We4HR��\,$+��4&=*��	�
wQ�8hE�۟F��� ���U伪 /�x�JsH�x����>Iu<��S{}��t�T��'��wd��8G��V2�E��Z̝��,��:9A��{��=�f1�g����>*}�/��"�|��:���:E����76���3Ez1��r��8�
�B1��rS�^��n�s�N����I�Z=�����=t��4�?��x?�Kx󭷮������h�):��>�&rn�=���/V���bw��.����t��33���5�u��3=�t~�k� ���MD��c���I��n��cps����6�J�D�y0�\d0����~I��b���IOӾ	�C�8�M���9���Źyܾ}��ܧ�\�[_��2��@�H1��$$�tY�e����%�j���^
��\��x��(�FC1��sKh�t�"/�����P�1ؼ�b�bv�<6��э�K H1=]�_(���wf�\	q�G�b�.�F��Y���q����;z�Y�w�qq�$Iz�uxuj�0S�	�j�wwG���ﾄ� B����an����iT�˸x�����5mIi:^4F4�
���K#k{(��22�o���)��!�/�4�Q�u����Kcxi��L0���+�'�C�d����� 8��2����e�7�����ܯ r���_���9��E�$u���/��	�;��S��}�l'�r�Pd~�Рtb6�L�L�+���x�/���v��'��m0��v�j���QR���@x�>4���1~���'��������>J��(Tt�e�ݫ)�=����㈗�fF��..��2�=��.x��:=$�E/���9u��T"^f��e��8�.(�b��u��X)N/�#\/�Yt>?���~���ǓO<���F��S�ykk��_����w�OZ%?�g����'Ly�b���^Q����gggmm�? S�c�ُ���,/�[���׿��?���($}$AK����)8i��<��f���ҽ����:h����x�*����rf��J������U��?�(���0­]��I��(���ob�v�3r)����݃F�r�� /A�Mc��ߙĸ�6��.^���(��X\\�b����"ɥ�p�f��+[ʗN/#[
��d�' �B��^y�PT�{���r z�����SH��1��^��^\�R�{�(������#�-^����Q�n�Ӎ�Lܩ,���=� _`)�8x�M�x�G�F��ˈD��/�"�ן���u�X�ų^-���I;N� vq��&�}�~�e8����,L�Vs�����*�g�%
��蘾P��3�U�x��	)�!�Ͳ��L`=>�G<
�<R�Y�|a_�,�� /��ޞ|�����ߑ��L(r$%l�7y.^�px^����7��H����_��}� ��(q3�+����x��f�?'��X[�����!�R2r��T��1�\���^!�^�����Wg�
h�Ia��}����3$Wx��Q��u�ެd�6`i<��0�cDH�J�z!��t�&��uT����j�k�>�C�|+����5�xPxy�x�I�Y�c�C$���@�Gl�3/�����Ø%�����2;��ǈ��4F���W�&�vssSX�L�3���?.���/���S��?�t:�����淣Q|�C@a ����?��B�$�GzX���0�c��7H������8R��P<>��2s����?�Ͽ�7>��uTr1�~Ѱ���,J���p1fٳ�y�;���6�A�d���U�_��č0���斐6��]�
���&��U��� �F{0�{��iD�Cx��D�~QjA2�� o�{�F���N�;�U*���*�¥#�޻���#����P/ձ����_}O?�4F~���3W����BY��)fޘg����Ű�V#�x	����K#z��Pȹ�=I���/��(}�g�n���dw~cz~��{r�H��p���8竈>�� A�����?�x�O��ڗ�^�g�ɳ%&��Se���	���LO������D���9̽1?�b-�\���l'�[��9G���s�T3Y�x�e��L�1�6���@1�#N���pO�I��#6U�
�\�܆I`+L0D���}W�d��N�X�T��!��o�w_� �?�b�0ƽ�)8��0����r���K�=?�HF�\���$�#���u�u���s �o��\+��c*�*G�����U�g=� ��x����[�ig!��C�A�*F�+i��?��"^�!�>^��ϔ��:2� Q�G�t���*\�N���;��@���������X����р#^ac��ד�"M5��b�7���J�X����\G1{�����5�,hN���
rt�N�*�A^ׅ�0���P�w{{[�f���=Nv�K/�$
u�\���?��G��_�Շ��o��Ɉ�� 3a�f��h�{�N�*��}�m...~�����پ� �o�z���������x��'�,��GN$���Π\�����fS�­����ܽ��A}'���.\� �i��3�L�S�ȓ�x��uăo �n�������SG����~��9ʾ*�:�[PĽ��V#�����'���@��ԏ�������V�������3��/_@m��wxY��EjS�6�e{�eHJtg��R*���#ℽ;���[���s]L�0ռ�>�c�Y����*�p^�>���;l�q#x0K�KI5�f�#*T1�+�j�y��z��^}��.�Uk_ƥu���7���OL�m�#lo�`���z�M��|ו��1[G���s�sR{&��b�k�s�A_'��`25���Ff�`��K#��xً;�����(�+%�J�/(��(�Ij��
I�Ӵth&KQ�,W�K��b	����p��`_�\�=�o#���-��9��u؀W~3�?���Ϡ��T�0f���aJK[�B��$�zC^���}9�j�,o��/��6n#^��-�e|��#lm��a��k<~�,�����ӟ�>K(��(�g�UY�M��� n7bu�Z�?z��-8[��Q�y��9l���1��9�άI��#m�������B[�<�:F�(���"�����/J�c���L��g*�X	�\,�9Q�S͡ .��稆fE^������@L_{�����˿$�dʌr���2����xQm�¹s�L��p�֍`uu�KW�\��`�,7��~ �������W���?�m{��/��0�Q/�P����*XZ�����y�dw��1�[�q�1p���:�/����(�8�X� �"�=J�B~��{8�6qss���4�������TmY��<ߌcc�4���G�M�G�*k�	�����b��6v�n������"ί�Ƿ��,~��� t"�]���tn��%���˔!�����x>*���iM8��)�D�L�	�]����(�RA_<뙹y���V<��T��摤�k�E��n�OVoF�
ĞT��1��Q���{JC�o ���f�Y8ޱ��e���.}�.}3�K�f�uLrkw�+�朙R��<㐼�`w� ��;x��wP�
4�<�f�2֎�|f��j&sY� RM����^���/�UZBF�1�(�$H�]�婢BD��Z)��/��Ȣf^,j$̱���6pW�O��wQ�0�Tsx���m��68�~�0���Y�ʟ��◰v�Ө��jU$ӯ�Ӱ�)`&`�Fr�Q�h5�9��ݝ��̖�|�������U�V��'���̨�#�VFV��m�6[�/���ڝ�x��b>���˭j�����@ۮ4NA;�`���C�A����ֻ(�!�M
{(O�x��<��_�f��<}�[��6� �8�疤��t3�k�L�3�%����/!TG$Hr�FN�=�V��U�k�(�=�q��N��\>/ j#^΂&��K���5\R���"�A��k�/�����]�cR+>��P�����(���z1����d{�BIx%�~Gdi/^���~��?� ���&?�\�{��t�p&�����B�Z__o�_�������~���������RC���5�x��V��2���`�y��m��#�7���ll��#W?D���;u�3��4�d��z��>���zo�hx��ou�/}��e<��[���������u�Vg��[�b�� 3�Ut;�7��s���ml����^���������)~��h����1�4#7k��1��ޖT�;��sRߡ!,���=�����]�\e�25 R����7�z$�M�ј����5[���yn���قh��I�uw_k�E�銨W���pH<g�z�o�+�E�*��)�x��6��\��ױ��Y�/\�a�2L<�Ɉ�>�T��>U
�G�Gy��]���<JŢ�|	���]��}��k��9��c9�����KXϾ>�z�jzxmK�(Tɼ`v�P�����CģHX��2Ph��kB�g7u�DGG��������|�MU�(0�N���ڨ��'�1rv��[p��*=B�l��k��Py3��������*����8&��� t��?G�ͱ%��ڭ6�>�aMǡV-��C*�²��%��$�v�C!\���Z����H��u<n�a�}�4����{qw���HKOe)%�Ϲ�.�U��9������K��x�4��pk^� hc�?�q�\��C��>
^n��Y�'1��)T90��#����� ����g��fڗ��s\�!�8�t3,O�[�%��kqh�����>��6
�2�gg䞵�$�,3X"g���3�C�+�-9T�y�V�#����u\�z� �X$��T8������B:X�>�����/����������K�� v�#�͜ԃ��������7���;��L�a���4S������K��{�\(�]o�_���/F��e��Qc��$���f��+�o��§7��q��m��    IDAT�=黛Y��r���5��.�v���(���h�'}�eT�^�꣗�p�l��4_�W�Q��\���M�Ns��8h��ft���(��0����OE�߅w7�ߨ`������a��=A�^F��c�㿜6o��νm���X^X�ׯ|�+x��������ņ܌�"�簵���` l~qAnP	�!or�/0����C4�5 $㸋�woyd���83?'�f�nu?���J)hw���V>8�����rϗ}L�TP�P����E���$i��.�r�;�7�x=�i��wI0��+�~˟���e�3�XA����,�d���'L��8@�n�n{;��H[��55N"@0m.Qx�'��*�4�����-�x��R�Z&�oA7Ǚ��!v���g�x����}�KL���L�Jz��KGIF�%����%	ԩl�Q��������=A��#`땎��v��(WS��8h_@��8ӏ���ǑzU��r0-!*I�b�I!��4pr�
�CD��`(�O�6�&��=3��K��/L]�}��8�i*ue��=;��z�zS�w�3-E�1U����2f#儂�%���2T^�~X���?��/��]��' � �!�j����G��
¤�N1_�N����ի�M7��2N�2�"�9�E�*�E� �"
9��d�Q4�gk�d���FꕊN�b���͵ȵck�:���ZU"Y[��9�9	��9�S՚���9q=Y�\�G'G"��#ԧ�z��;��B�����$��u��~I��\�y�C�h��&�*�o}������q?���x�e���\}��W�8qݏ�0�-���޻7�u�D�T#�0U�/,tWWVzΝo-/�������z�\oЙ������n��*���b� 8�6�~WH.Ӌ+��f�4w�q�V��B�x=o{�������×�H��/#-Wx/D��.�V�gt�{/����5Oc\�g?�7�/4x�թ�IV'�!�V������(1]�3�pw�o��+/����4y�Q|�Ͼ�O>�	�dV�/aa��U�%�w��}t{=I͒��z��W3uT��MKq��Դ4���<�)�T�sIagLux	Z��`��u�r�{����Q�E��bz����1�D��P�P���PvP� D���I����� �o�8u nEN�����.m�2V?�z㲈���p�3bo���s�<h�٧Is�2e��<>��4��F�DEY��p�x)g)ѓ��&�q:*l)�"�^�7�>�Ѱ�sI�����K��ib�(r��;�X�rEU�M����}���BNK�.\/B<�y��`N���T^q��B������}��B哨U���Ǒ����d���ȕ�n��>q��� S<$�eE�F�#9fz�]��]��GN��:t<�����ű��c��'�O���D�g4K��66^ِl��0���8X� N�Cs�ԍG"cI�E�!Y�ܶ�r�"�2H^r#�N�4�sy�?��Ǝ�c��C ���Y��`�0���:"o��֦0�F�D�H������r�TjzOyJX�O�!1,��d�� �AT;�J���J}��O�g���42���Le��$���(�g0�|sS�Uz��7k�A��W�L7���9���	ח���A�q�l�uZ��&�&?��t:���b?��_��g>�aa6�Ƣ������֍w~��C��'���SʣQO6'���Y��a���O�.��Yȣ�k�_�C�|�e<zy�~
?�"t1��L/�X�cya���'x��ȵ��k�;�h����ױ|}n�NՂ\�l}w��`+�$c������Z�<�Q�?� ����U�^M�{���c>��C�~�A�� #Ô[��r���$<��믾�j�"-�z�[ظ�9��95hIIB�bE��oo�ddɴ/a�"M����V��P(<*����ޮD:a��`�L� 8i�ľнC�1�aS���Ĩ�+��
>���~���8<>D���;A��B�q�p(��u�{'Do`��3X9��(O�����U0a�r�
�t`�F�D{e-�Ұ�� N	����^dc��)?�.��e���N݊�4�X���������3'q�2*f��K c����/)E��yd֫5JK�Z{��J*��	�N$z���n��-T}��X���9�!���T���O�/6 ?��ij2nCIȪw	E���Ԍ\�wC�I7#QP�# ��{hLϠ?�HR�U~E�{�l�<��7�GP<D�̑�2�*ck���~WD61r-�3��|�I#�ֵ��@�sDp�}�����(���yf2O��r$��n,�)��aș�Lӟ��(�:�J=�JjW��yƇ�Ea8��ΣR�BDau7�0J��N�fW��T�5�����K���C<�c�iZY��SU�|l�{����'S��%�@$;�$���$ŋé[�D��n����n*pK������p�e��+h�O�:aWA���g�Q�ő� ��N�e+��I���r�>�Ao����/}�s���̜�X���;��j��������$��SO���q�#v KZ�|�ۗ�t4�x���u�.��O� wn� _x�Q��6
� �P��
�)xN+��p�C����(��"�w�H���v��.�zԓM��I��A��я��vu�nas����A���/!�/�ᇿ�eXgv�T���#ؒ�RE��oF�$HQ)P 8>hbks��4�S������s�`���Jv�Dd��
l�l됄(��@��x�W�fs�#�>��H ����L���tt�o��	�H��������
A�����5Fu��hً�av�� �s���C�s� -T�"Tg�pˇ@)F�-��v�8�,Sb�־�ru���l�X���&=�qz�6RR~*�(Q}�lYF�2��ω�_"AN"��D\<�X�&Sz<V:65����3mM�����x��#�e�$k|�haM�#�ث#f�&�U��#��g:�I����y�!8윬�4�2U8
p�i�� r[���b#�~~�~R��;N�Y8�*.�=�JmN./�lciv!娈R�*�f1��<���=8I���&�Dk���:5��(>�e���4[�f��-���� �f[~�^�����y'۶��`��vv�p��Hm��S����:9F����Wk���'Az��0u;���@�,\�N�����I���������R9/�`i�A^��L���X�P�JP(�(UjHӒd��""�-X98>S��A��06:����$le:�<�t�R�u����k�JBc%��-u�m��֯���\m3����2�\���a6�틠F��A0Q�U��'�>aϗ��g>�Y$)k�O���@B����%���fZ��(�sx���j?��<~aq��_1��Xn�#�U���?����.������?/c����EK :�H�ɨ��a3&����x�-���ve���o|��y�<��%ԓ
	k>t;=8^	�s8���?B����p~�C�q��t�+��zuN�A��@!:���)$e*�qa��a��o"Ώ��������%ll|�<=���>֧|����^o�r�G4���9"��u��&�{���z�����f�rT.`aiA�������]���:$��yM��9�M�t�	4|O�`��'�a����}| �fkwt h['�T��;�; <:A	��K��lw��h�]�̑Y;��0�U�=F;:�ܪ��E��t�G�9��G�+(���/��XG�fK''�D�?@ЏEĞ�U�TA.�a�)���.�������J��ȉ�mӠL��-p�=	<T�Rg��5�˵2�����AMV*����']��#��XaJؗH�S�"1�<5� �:qF�J�YӬt$+�Z��=��P���D���N���D��?Dc� �8��"�9�؎p�-"jX\��be�bIf�r?nݼ�h�,@�[��J�+E@�}�'�e}H���x4�O�ϖ�(WU�Xf��E��c;=*W%�V9���J%[<���qS��7_�}*x�$/F�d�K]�' 1�����kZ%��k���|G���}֘KEDi$�ϒ�a�SIA�W�ȇIp�<3�M9�P.`���5�2	�#����2&�[���nQ$��ŵ�{�3�q͎�����fFd��x���?�dK�9 YY?+����� A��f;U�J:`��?�k	�t��(�eAHu�/�I�6GLj�Du��� ʬn��%�4��}�֧�-�����Sk��}(Z�>^�ݻ��W���������4��[f����7ޓ��� �|(�(�$Ȼn���^�:S�1^x���{8?_A5�Ï�"C���� X���b�b:�0<؁�����i��)̬o`��81�u�x��p �Q�W�y],^�������ƝcL7>�N��{��\���O�P�0��e$��`���{!>�L�1`�#��E���dr����x������ۨ�a���~I�d2u)?�:9���$N١qdڎ7,of�����0wUp%���`N:B��C���Pp<�lͽ=�$o�Pb�E��|�Qg=�G�m)�P�/���B� NC4�M4'hM,�50���F�Q����!���,�V�@���T��p�l��u�5���z�1�`{�4�6�]Q�a�+�ٴ�8,���9X2�o7�������.��X�p	�����r=p�3��F�C�/;�Ϲ�/-'�D��N�.!�r_"�.��H��Zo��C���5�Z&��#G�u}�`�$���z}�yFP�����)Q�>�q	pr����AI�`��L�C��	����D���5r:,��k#4��h�6�#�V1k��1�,#�HX�-I�R���t��s���u呶W赵J'�ڴ�����%�O&��>��R�c��r�����1�ڗ�*#���z��\�H���8v�C��fF��"9R�ˑ��Ȣmک^�줯�o�S*�!-E"6���$�ڶ,��H�
�ک�*��6�wÄe+O��	���)ݞ��^(�?�z� A�vB� �YݝΉD��t;X���׾�|ᩧ���+���2D�+ީ���{��=���<������'153�����!IP6���Y�9.��(i��p�wp~~	S���<���WZ��'������P���."&�w\���0
z���AZ�a��:.]�����{�P(�9�¯W�O���^.�d��@�so���J�!籼�0j�y�.+8>�`��H�M�D?�|,��
��=��J��Y��N�����8w�޻qK絲vX,�GC����5��ӑD�DǜkZ,��I��ݻw��k�����5�Sq�o�H�/"�_�҉щ��(���6�N�N��
��"�5ʒ�lu%:`���� `���8t��n8D;n���f�kpK#��A���$�I�����j�r���0��aͣ6��W�P���8�y�0dj�7��<.��x"HoH��v���l+*�j��V�����5^�n	VLAK�b�MC�ԈQ4c�L��{.��EN�"x�dn+��,Ј���@#fv��+����z!��� �^�G���n_���i�
�}*C�[�`0�4��F�Mi�	
L��c �۴�ީ��/��K-��b���En�s�m;��O���T+Y[l�"������v!�����-ۙ�bF��T+�e�Ӷ���O P�����rq�)��0eKRW"�_��ٹL���G�gM�}��jŬV���i�Q�ZɘQc��J� 8�+��g�!�IO�\W�����V*>�,���g�����aMV~���a8�k�5�P8�(k�6�5]>8���@�)�k��R���(��}��E��gK���D����_�g?�ߺta�w��1��rs/�͝�O�k����%<��Ϣ/}f�0����s�Dl��MC%���{���.-��Q���p�Bn4D���`�Q "D��)c*WG=_���st�^�D�F�4�eL-/����lwo�'7S/"7]����*��M�e���wol#_��������f%�Y�M����Ξ�	�F��Y��P%)�>UA��ł����B� #�b�����Ćx�ݛo�)S���Ψi,ތ���dŔ�:I7	�R#]���TCCD#@�$<$4���FR��(��Ȗ��U����d�b���#S'D�N6�\
��)g��8V�6��%�.+�FN��r-h�9x@��w�ɔ$�σD
�zb�u������&ƈQ�i��[N�A�Yf�.�k�K��G4�4"_���8B��kjy\�#�]R���j�N���e� ���Z̢9M3�2M�&�̆YO�+Y�iݖ���1�H�|bE`MZOE[�J�)a��5FG�H@�,+����������x:%S)��~�� 9W�<$�ѧL��e�s�Ly��������s�kŴ�c֏�����4׀y���Թ�3�2J$�s���ml���n�`D.�m��9���PF���&k��u3�38��.봒�����>�����)qb�p�Z[f-X�GN��2�$��ͣ��q��*��,�%�|)���f�: �w��mK�n7���.\�X[ ��j�ncfj����]��_]�|�C1��#�p���_��?�ʿ�]Z��x)gG��?�H�F��{^�L�A����z�V�a�RC��ī���a���tI�/Q/�i�p�^n���V�)'�#�g��r!R�F�@aQ�g�W��>�J#?� �!m��rS5)x��nρ_�F/o�j�&��ސ��(�XV�W�cgDT,�0tP+0�uA�G��F���L�B)޲Q]"�Q����.}�њ�!���Wք%�r���a�jk��k�F�Fxd����S�����2}�T�Z,�A�!E(Z�Xz�y^xň?$`W�[>�)��GL�H-`!P�Hz�i-���/�Y̵yXeCp�
�j� e*�:A�SZ�xy>���J�aWL�9��Y?���[X�W4�]��d�v6ұPzQ��J
���w�-��S� ݮ����$�%-�k!iZ�r�˕5@�;\��N+`�u�x�WE"W�o�O�vЈu��f��=�}e�g�fJܲ�-@�χ�V�O��'ۆx[ڶ+<������D>�/u�D��[��u��*]@�9֕y_��JWz���5�lu�c��5��=.9{�}�e�����ɽ�N�y�d�~h�đ4�,mF��p�~���v)��$P��lt�lT>�I"	���IQ_���$L�a����1]��W^���������0��O�?>^ ���w��������~������P����7w��/�+i� l�H�4��K/`�1/�ATP��/��:¹�E�I0rF*�����L��Pt��.����9OU%//_�����8�o#7A�� �h�lT�Y$$���H����$�H�	r�7H�a�mD���uȔ��Lʓ����`r��	;��D&ܮ&`��״*{l���<�	�*�0�/Km��ZvhX��
��Z"��3�K�# ˔#���*"�]�1vܶ9аUBX\'!��$`H�!3� �/���	�6 L�B"F�AMo���nI�Ka�fڀ�N��L}�X��SGC��2�T��QR�uʹh����4r��ŘJ��%���a�:�^�O��ipx%r�u� 	��_���O��`���#1�:`�92Z�k���%0dfB���3\���l"Q��_�I�1���̯`]��^F�&0�i�����,���SN]&� ��\���� l��n�Qi��P$�q
R̆�T0�+��kB�<�\Iñq���d�m�H��1�N��=Y�� /6�|�:�"4�^���}�m	y^�x�y��vfSϕ��l�)�5^�]�0���5>�|��\�~E�/�k���;"���[o�����te����)��ɽ�a8ȿ�wvv�oon���tV���|~Mҗ�l�%��i��H���:x��P/V���7����^{�u��._����Y,�.�P�bH���A�P�T����(�2-��MT��1a��1	34�������    IDAT�U.dD�`���R�6s<�B�Q�0�id�7ob�z@#��&"&���������Q�M�G�˩��4c����&Z�[��JN��@6�C'��5,5��"%�JBp�1ӡ5�%�#'�h:MRt�2v� c�F��� X@��F#s1��u�+���o�JzV�L�i'!�Zթ$b�j[�0��#�cv�2��Q�7�+*B�$b�UHB���q�`�Ev���f@;�UC�1��k�5ȧ�6���S�DY\��<q>���2�h<�e�;����cT�h[��-�55z��%�I��J8��	�������lD�SqtL�#��=oR6��,�d���v���,�V���\�m�f�����dB$+�C�o���'���qG	���{:�l�T�׆=����� [�=����k�,�Z�)[�,�)�N��-�Y�l�MoCJS�7M���'�k_>�O��}�
ܿ{�33�{�҅�l�>�q��g��w��f��Cj��R!��@T�H��n���i"����s��#�Z.Ґ��s�vQ���$��RĬ��DE�=%���bm����7��uK����^?��M�7ĸ�h!����I ��N�B i?ǈγ�P��_�_{��\xf�\$�8J���S+��"ӈ	��
cО��Kc�a���8k˄�9�z�;!��pf�SOMT�Ԫ:tv���kӯ�m�N�Fw��j@T0�FY�Ό�x ���\ �v��q���@ 2`'.�7Ҙ�DYR������e6��u9i�1����댦�f�s6�,������D����}�3��$5훔�È^���gk����j���Ѡ>E>�7��U�/I����:Hⴐ7O���F�	����86j{P�i��8ⷄ�qZ�83��1��F��K�����!̚8Oʀ�:BBHJ��Y�<R����hێ��;�f�rn�u�	�Neulk�����<�2�ca��L�l�F���f���s4����7�ŀ����vdğf�]���mN�`j���=#�Z�q*`1�}�Gt����aBmq��[*�񵍵_y�����ڇx_�������G�\��I^�$����Mꎁ�ј�~,3�g�I�����
y��=I���sBRĞ��Nnʒ���i?a�7Q��\؏)�T�.�yհ��71���.ۦ%S[�1�ɍ�e4D�c���$:�U"CX�*
Zg���f����ذ5}�lT�M/��¬ͤ��o�5B���F/�����pSS���F�Q���66`�5C�;#V;Q��$�ZCTC�5T������٫�RԤ��>0u..Ĥ��29[��uN"ӷl�3�<e��L�����FR��ݳ�=Y#$����&}�=��mۄ�+c�X�0��#0%�%n�(�C"`��I�����E_X�#Ge�����	���p\�~��+�@�	ةؔ^~��9��d?g_��]�=ȁ���@wx�������LF��K%��X(��T	dR��4��P�s�D�Yj0���kl#~{�ς�u�Q�]7ܖM#g�Nv}��Z��{ǈ���+a�Y�%Y����IS#���#[�}�l)���>& ���(�t��-;/<te�S?m ������׾�����C�����[M8ԙ��縬p*�NFGw��Ŧ�����F��ϔ3!�i�`��Me۬SUr%��C2�MO"E$H֠ns0�x5M����q%�~J}�S�r]�+PT_?�����h%���$ꈥVLs�7�����f�Q@���j*V�o�r$�����T\���ޓ5�h�e����YS�uF
AL��)�ͤD%�v��T[r$�LE�_�+Xo�t�g�A$��O�]H�T+�U�H�%Ӭ4��?U�zM=K�^��H�4Q�!Id�1�r��j��NG'j���gӁY�x�.wH�.�y�M���JO�DZz����*$B�IP�W-`��1���v��&,�<�Q^'�8�1���t4�JL7�!��X4���\o��G���ᜲ�K��Md���O��c�7{�d%"3����b�6�,�xdץ=/�h�Fx���N/N+�S���Me�ulr�e^#]WpSޡ3��O������:Y��-{�-��}&7#됱�F��5��j��ө�	3[Jf��-!U�����&SY:L�8KD5��\Of��͞'SN��t��f��'>!ٻ�3 �W�JDa���W7���3�o|�߸��WW1�b��+���,`�x�7��P>��5%�!)�M�l�ѻ���Iհ]g�91 ���u�ry��4���5YT i�P�!�Jҩ&E�1h�r]��$ulHD���� �Ɯ-5|_ZHt�-A��i|�Pf��k���Í�k$d+
p��?�D�B^�	~Ph������e�J;��$�Sc���߲}hl݋��v�7�"�S.OSx$Mi}��$ړԶ�e����(��!�3k��g����i�:�6b9^�Z�4ǩf�#MJ:L���Y��)�jR��h��ؑ��~���gE[�Q������Z�<��,!D2� �R��~ �H]��P��N]�>\3�J�@�FĚH���<M]$i��.:A<����v�.H$�ߝ���ڙ,�M5�u ΍![q�J×�S�����S�#��Ҷ���Y0�v#J��3tp�Kf�h��}*iz�)2�+Ζp*�&�����~^��� �e%�˙�g)�'��06�d�L�i�IIN�E��Y��!��;�VIU`{�IYs��^�1�L�p���W`?~�:2!K������r�0F��c�=6�H���X��f���r~���K����Ǉ>����~�_l\��7Wέ`�e@��3�+RQ��o�x��E��\�ڰ.�ӣ.���� R���YZO����c#����z�+#5ڈ�b��L_kQ-��3�D�'{����C��ٔ��4Ȝ�-�^�&'[4;�YȶL$6�c�[�'ӎa&M�cY�r�I�2�O�T�[S�����K4;�oU���A�K�b�(G�����M� J���8E��4~�{��]aK�T6�l3a��qL"�o�X�iϥ��I���.h�#����޶+���%eʠ��;5�B3�QJ�J�ʺ6�l��Ð�d��Ah��k��dM�M�+���^��y�dQ`�r���3牘'�kDAd�L��n�l���q
;K��_J�m]�,h��*���F;b� {V�(f��~1
�EU����G�0�%���Y�&�d�����W���F�F��\�q�����ҵ�j�a�zŤP#N���5��ͦ�J���k`�-����(�k�% �|�Ym�J���)�I����̧d�l)���Q��t{���^<��P��h����z��ʟ}��6�^�Of��sДToxI��N�48V�LQ�>�v�$#!?u�t�%�3�7��8�˦�.�'	�*�gH=&�f���P��h�ɍ9�4O_Z��e��7��M��D�7�%Ai�8�۾n�_Ҽ"��!�<x�|H�e{W3iz_�
�V#qRX�D��ک��m�u)#&�(��F�B�~��ɘ�q�����:��͂#��Cj�&�GkF�A�AH2j�iŤXa�Ɏ��Sj�ڞe{oD�`�W:7�5%����k۶C�K�w$`cj��9�R�z�:=) !Αi��\��H%=?i��f<	T4b�N�f��T"\S��Կm��X��zڵy�YWڤ`�lq.��*���R3&�| dr����$$�kE9!.�r����V9+[_�smׂ�?i%�t�e��ʕ^�O���c3�"S��ڸu��P���n�T����排�a��	�tx��A�$��>$�.�J%V�+���2k��4�u-��~�ӟ�n�{)�#}�a���v6�6W^XX��)�ۉ��i?�������g��ڕ+��h`��~�$�]�Ŋ��&��燀���mh������Mkk)d+K���f��xT˳QL�N���)X����51�8�f��q*WR���ʦ$O7غ�z�޿��������9�Ƶ�5�b�i~aXA�J�d�L�xl�`�=0�  �ϊ��!� ����c<���{%�Qe�R��
O$�F5kC�IqR�Xڰ�W\���k��ĵ�P&YbU�9��;v,�I�~x�r���f�0L�e����ә����=��:1�k���H������w&���FƲ�35ahY��,��Fj��t5J��%ub�87�,{O�P�hi��c>�,��w	G�mϻɤ���j9 ��[�E#o��B�3��m�co��1�33���i�Օ�m�����|�0�Je��~Aցo�q�D��r���hLĴY��4�e����{x�'�79Q��F��-����f]^^��~��O��>��?��?^>���R	G'mT���)sMys&x���鞍x� �1��W��l��E�z�b�Ǟ�x)�H�DZ7�g�����{
�m_g�Eu�M�Y1�G��, eA��g��_��H�4	�A�k_�흎|����/+7(�*#�0�V&}-�3l�!�T��>u<�L�_�WY�bЄ�;i7�z�IK�a�Ξ�1���,�*@�@*���4�B�K����@�6k˴��qPD��L�M��f��H4/����^#�w���A ;���}�����e�O֏�/��0�v_��σ֨��c�7Ձ���W�V�1�P^���(����:Hh��5	I-���̽�k�5�'UG[?�R��k��<��6��-�0bV�Rfܴ�nF�f���U�@�3�A��1��r���ۢ�lץ���7�o���#8q��4�̈6����O|��!$���95�=��Lc���pa��ɕ���~R�����x���������Q�%����6p���5�%�6D�j�jo^E�E%�UB�x3���S�xٞ�~�7Ӂ��p&����)�̮
c���Ѓ����|��߬�9�3g��مi����'d��7�9��"l��D.��	�k�D.�Q'��r�ykȳ��$�"�[��Y���EL�D"�2��j�X��Sg?o�~�N�ݟS��]�Q9%#��ޤ�ib�SQ�"F*P�ȁ�
��h��m�h�N��T�6�>tjZx~�����r���A�@����̡͌���e/�=&�A�8i�k��x�.x��}"�7fxƺas3� ��p�0�2��HW���%N��&?#��@�kLA��5� uc��u���z�>k�]{M�U-�ĉ��l�G��X�C�l�q�0���ߦ���ص)���4�{��jΗ�2��K���4iu�5"�nmm��#�X�4�>�(q�r�c���3�^^^~���O��>�����/�������!��K+�F�/�ۈ�Z-�
�ʨ1ⵂ�x�8���� ���(�	2d%x-�9kl�^����8U�<{a��C�5 F2�� �y֐d�G�Y�y
3?`��F�A�ekV�0gA7�؈9�|�%�S`>fL��������|�V����t#�o�uL���uD�'�&3�G�D�lvĉ0}�V�?+�8v��N�Q�2�K���8{��5f��f�׏�$�$9��:�%��7�Pgd-�$24�f�G���R(�Tt8NQ��A�$��X�Mm#Ks0�}b��R�C#X[+��t��"MM]ײP��&�t��Ǫ���$�T��0'9[b�|��k���jń@05<I���ʒ�=f{��T$��8M/�*��}ٖ�mP�ҁp(ޣן�mD���T����T���3#e�c��تR���L=vL1dQ�9��M�e�q��HM�}9���>��l�5^��O����?�I����z��ދ���++������|N�F���r���ͦ���bgX::�SسF�����$LM�;��Y��t��xYW� �<(�|P���2�g�;��V��e_���cl��>h����������8��SY��n�Ԙ��� �R�c�w:�������ˤ�&�ղ�M�R�Q��l��=����w)Qh��k����`������;&�'�1�h<�����흶׊�|%����$��o�i��ڰ�lȐ��҆9
�T�rl��JX2U���^���xd�Y�Щ@:I��<�e��(��G6�y��ۿ��'�;RD��`)3��`��i�]�WR��5u��,H��S%�[ވ�����𘎺h�ۛ�f�x���6
�rލs&��c��U2t|�(��b����a������J�+�ޒl#o�v���ܭ�u���3#br`h��rޱD�T�ⵡ�ۻ2,j�~����Ύ��jF��lU�|t[�q�;7=��kkk�~�'�sz�}�Ņ�������6�W$R啘"�
��\�i&xE�� �ޔ�G�3-Vِ`h�8�X��(=�dX��m�9���W���bF�=��zT� xf���X�X�wt����9�������')@��-pL"�SD�A�����X������_6�2��6R]�qː�u��t6ړAL�O{�4�ۤ�h������CM���J��,��?kF�e�2������@���<F���o-xg{B�{��N�IA۶3[��^[��tU�?�+f'�d5�e���LfN�95���b:�^PL����Y�]09��}f�����;+cUǜ=���?e���8�L�[�]6 <mJ��ȷ��<����Y�2���N�@�s�]����y��i���� � U��6�i=�	����iK��Q��u�-��}��"�}����##������4�:8_*bzzF��A%|�8I
�L�Q�A_��ҥK��e7�N�p��N�ccc�������=�>������˿z���R��M0!<�+�s�6�'�f�" ���Lb����Q��$��M�̺�76O8ӣT��|��٦A�1�eRM6�*<�S,c<M��M�e���f�����.;'�o��ٖ��gSj��$�U�HI��^DLۊu#��Z���'o����X��R& ���˴m;|"i��q6j?����g���4�a�-���P�CTČ���M����; Y����e[@?��v��̡=��5PQ�")MF�v�E�;�~v��u�t���p[b�|��D�<�.dJ�g�Т�����$d�Fq���Mۖ�1�L�qP��k��v߳�r��v-Fq(u}�#כ�3��wM��g��Q�"�&�#��IYD��<O�� ��n� ���шT��Beqƥ�>qJ��+'5�>��汓��v�O��mI]�$���@"�*�{,�e���a�m�	mEy�cq~���6�O���n�BA���0�;�u��(��m\����I�F�^g��9�muuKKKB��m-��>굊��g�ko���?z� ����=�~��翾v�򗎻�1����E#`h����^'����4z%�ں�ވjP�b�����b�X�q}�A�L/��I��F 3� %iB;���yL�P���Y�6��5ʧ������k�o�D �L!D����r\c֔��'�@ȺO&x�����̀rkܬÐ?;�����&��M���G���d�5��%�5 nARR�&�;K���ma����-��5]��4c��&r~\6��w��@��D�q��Ԏ�F2�x��6��p����?�VM�Umg[�d�M�Ħ�-��v4���o��\�H����y�L�S:���,Y�=�reE��(߳b���HFY�S$7��$JK�X,([:�����H?},���}�"%�)!�q��:
�
癣�>�o�&�4'S:ъL���O�71;����}��%�#\+�'@>���J�����8�0{{������|q4!�Y�_�S������k�9�fp��8�]�N����L3a�/|�i<��'������f"_�x������(}�w�2��A	����R*��_��;?���~��C��|�{�Z�v�)���K�x��:�q��x�Nd#^+�A�e*FR-ƨ��;1�d��K�*	Y-�I�z��g��Ƈ7�����l��Yi?{�dAj�IiV�J3�.�Y-�,����^@Kǂ����e-#�`I,�vd[�<��ٿ��l$v�������M��uex�Ti&ҵ_W%�q9v�5֡��5:n�    IDAT���Q��=�-�� ��ڪ����s�x�q�&�<�T�Q��5B������"*�f��ݙ�J������O֖e�f3���E���]�5>v|d(�e~F�D@ʞS� �u��]����pc2+ڨ��^Չ��)��u$YS$�HM�Hwg�B���������# ͈sȩ_�hLL�Dx�b��u�l�.�U��P
MH-���ܢ�o�G�܎0
�3MT�.�2�W���Qo����������*�Y��ts9ь�9��}�D�R	�à�Z�l&�5d��5�Rǥm	#������[9n��̔���ӹ`�J���3��: ~���� o��U�1O	]��w�1�����xa5S@�Xȡy��M��������{Wz^g���s�97Bw��9�lf��(K��G���z���r���*��S3;S���뤱d�eQY"%&�Q$��sD#�ܜ��y/n7��n�_���.4�{�������<�9���/��>������gڻ���I�,^��\��+&�����Jn����\Qjۢ�j�F��*��t�"^P��L���vF�U��aJ�y�n���#��������i5���{����m�v~���h�ߙyV3^�UU��o��R�R���M�d��5g�j�i���m�RQJ]UU��
�V����Y�z�ێMB�����_I��~>T_��f�V\1S�fT���s��}zQ�����fW�>���/���.T3�j ��������kQk��T[ժ��TK��C���ۢ�*5_�Ū��j֯(`���T2pY�mE�
vx!�Za5���rH=tۦ�Zk��h�N���Vk�MŪi^��=�(Н�S����ܕ�6U
����\���U�Xe��X��~  &ϩf��	d�V�ʸɪP��5oG�b����yrog�iP2)Loғ/�1[͊S}��u�T�L^g ]�+Z"T�)�H�+�(�F�E�]Ơ����Ӎ�M�ڠ'�Ia��Ȋo�xʋ۞j	�zeW2r?�z��i+A��k۽�"���"��Lb�քս���F���f�+�ݽo�d2�~�Q�x�o����v8���W�f�����*��!�HO���?��
���u��ܥ��ڻ�J�+�f�/��ITD���ޝ5���m�i��Z5���yQ�mG��*�ꨐ��ϒM�H%��搈sg�l�A\ʝu�����J}e��o;��!����k{d���F��I3�<�V[�v�p���A*}}£U���3ם_����ɪ�y�����?�Y+tc�'`G�Z���l�Yx+5ӊ��үx�}���
5]Vn�6�JT�Tܹ+��s�m���촺~����
*sWw���#��_�w�Y��iQ��v��*u���L����'�����g�6���dNj-���P{)�Kjի��a�Ϫ�U�r����.  塚��@,|keĄU�LV W�.���s�4����Hڈ������Ug��T�bd�2x������O+��{�_�6+ RT$˫�T�C�`M���5�ߓ�����e�D�,�+�v�\	Rt䳅� IեKbE���-�����ihM�<��|)Si
MVR%-Yޢ��JN�2a��Z�)U��sZ�9D�ԹSLF�3�(H�c:
J�"-D�-p0�m�&�Ţ�ڐ�@A|���H�V��&Ke���H$���ו��<&���J��L�+�JEv184�3�<˾��dr��Ǫ��L^�Ū�f��
{#�B>-ٺ�|:I)����ݟ�E��qz�=s������"��&S��xŗ�^��'H[X/7|.�!��P(�(d2�2iҩ�X�D<J&���0� w�f ��=�;_9�u���J-�z�*�wY�Y�����:�[�O�l�j��z��%�:���ȣRC���U����r����^���ݧ��*x�c'��3s�v����{�����L���j=U*S5��(S՜�{S]����듬�p�dTfy/��Q����E0*�R}��X����m�7�b@PqT�햑��U�B�V2S��ۥ�*e/aDe4Fx� [��˴+�W�j�Q���2��ba��X���x�0���&�*W�2�X@B�X2O�2��"���7��_��/V��{uR�⥽N��Q���H�mA�2�������*��{,��,�*&���^:X�R�C�����x;��\>��������Xk]��^�גL�_@����U9A���w��L&��2�ER�$y�h�tV=e}I}�$�=�9�l%2�����k��eF+�P�P(F.-���->�YɼM�l1�Nl}�R.�t�LF䋀3����l����ڎ����rb�ۈ��LLL��j����Q���{������KL��+-K>[�xe_d3��:o��8N߮]�!��8�(fW	�Ԅ�lN�rH���L&�V�R�Q��l2N.�~ax��O���/z�z�}���K]}}���2^�^�j���%J�I��u��f�+C귝bd�KR�$b1R��h�T<��eD`�L����m*��ZV�A��J�3˽��(��̝U����
����^��[�O��T��?gkW�)ܾ>��Td��S���F�
����I���*pU�^�y���a��W�|d8}Uxv?�Tc� ���fJ���c��_KdEE��Im���ު��
NTG��� ��c��Y��n���T�V��۞szO�^�TJ�m��0ʽ��v���"v̀d9T�تx���W2�
�^�6�K֣ƽɞ�v:�w8Ȉ;�[)��sw���'�R ���lSf���g���V�Ѳ֨��e���%=���բH��2�G�>�
X$,d��(�|�re�Z�tU@��r�+nO*2l��U�@������jKLu�J�&�q�s5��ڥ^158WZvtZ���M@E �QL��'�El�
�7��ˇ��o�6Uj�i�:�<nJ�<��d.�Fl��6�֦��9��a��w�3ۙ_�3�fla���L}W?Z������[���K���RE
Y=�`+e�4�w�w�X�{���,�d�\:ECM ��@��b�� o����G]>���8zk�����r�����on�Z�C=�T�n�G#7�]��W_����ӊ�\�`Ǡ��'�bh�n;ʁ�UЪ9��u���'�����=+�q^��J&#�N�d���~Q �e}܇x�;s�r׮�a�vwR͒��G��+�Z����@f��*�э5^{�e�B�(qEY@H%��-�m7�J=W���e����nX�v��/kՋUfu�WjʊFV�8�J4)Y�v#�d"y9ԶM
���j_�������P����u����$�����x�]���%W�Z8���� ���VT���ZU�1����VN���2Y'�D�(M�UڍT.�$چ���;%n��m�CT:"U�R.�YI�W�0�87Ȓ�Ц%iӒ�(J�o��E�}��)���g�n*"@���a{"M�����=�xT��* Vۤ�\�=���le�+5���� ��E�&Rǉ�R�j�jƩ�6��ݏ*&0jm峴�+��k��%��7�O�P�!���6��d(��DFZ��R�"�����LAoQY[�,�I=�D�x8M&Y�XZZ�	Y��B�l"B6���V�\1���e*���wj�d1������ۭ �l6�ڡdSf�E��ttt��zp�޾}���~��ъ��lR �v�)�3l���ϖh����؀�����B��g���]X�T�����:�~��N������i�r�QƇzp8-���fj~���Y��8%s���,>�m��<^.ݙcn#��|�pV������J]K'�����Dh=9=[k)L�ʘ8t�8#��𵿧ߢ�N^Y���U�����o�����j����խ5���>���466���/����*�X��Ǐ�^�@MP���|p��g�q��)V���	S"���Re{�)���������+&DX�{=��^IB^���%	�3R�Ƶ~�*����v=��
���u��ܥ�W�[[�H����_�d����r���f	�No�`+�"�T�o<�5�W�ن�F���V�	U�ڮ���0�Lhre�Yq�*S2ŦŬ�a2Yd<�:r��� �E�h0Q���*KF�V֖:CEQ].fT֛ՙ(���rR�j���L"��(AAtv
�#jT��Ѡ%�I�����p.$��g�N��dґ+f0�*��B���k;Ӻ��-՚	�T��y�-�X\r؛�&��Dg�Ld)�E�Ӧ'��b2�0uʐD@Ȣ5P�y6�UԢ�܂ ���Ii�l6��$E]Zf�SC��T���j�l�Q O����S�HTb!����@��R�V��j��E+ڢ]^K&�%Z�Q������I���BM1��K�s����Z��.�U�+��lUԦXK6*�j=1�z�YF�	��S�]8���6	4� S�[�w��z^��)�T��ׁ�n����2�4[k��Y�ep��,���z�<"�S��d�zq�m��iL�b�խu
�"F����Z3E�/f6CInߜav����CM����nʙ2��3�g)Ɗh��F47���Ћ�eR�S�S[�m&,F^���!*W���H+Z�Dkw'�-�\vj���|�2�u�tw�(������ݸq�W_�1��>�]���yp�&'Ǚ�� �p��u��A�--����1v�:S7�[��\����c7��=8H__���"�.��\:��a&�`��y�_}���<�����b���V4�}�|����Kl����#%|�v�u�iho�#O}�/�+Lܞ������G�au�R�x��	���=ƿ�ÿ@��d��Ώ���Nʅ"{����?��_�-��,���w�f��~.;{�#�����/�Ne�������t*c�K.����x��wX]^��"��d|`:�B৞z�'������5Чd����V�be�*Et����������c�EHD��F��9���/��>������W����$�y�j�khP@�jWJU`llTe����p�i2Wzs)���_cn~�ň�b��Ia�j[¯�h[�aB�Eg�\��s�L�\S@'��HL$����N[�n�;�4F�z̉pB#�	�EQ:R� ��DAG���h0�`׉�R�#-���ԫ0�͛)�����hC)`��5��!��]^ ]Z���@��Z}�t>��f�l{W�������^�P�Dj<�P�D,���V��=�D2Gy}��*��.��jB.�T�I"���ɣ��it8tZ��ߙL*C��@:�#���wZ(b4	���2���H���-nesG�L^�'�ʐ�执u��g�yk�e%�)���DWsDV�������O�(��E�4��<��&VR����RӔ�Eo"�I��+YRKk+��Zf#~� \�p$��;{���P�Tq2�F�ܺy]emK���O�WJe��[�8�LL�i��ߋۢ�e5b�Ǧ3DV#,NΠMg�	�X��� ӳ3������tv���`����D��RؚL{؛�=2E��1&'C\_G_߅����Ǐ;Ѐ��a��<[3l.�����׸�[47u����ݥ�5Ej}�&����:�Z�$L���ק5i�����L[g�z���;w�����*T�˫(M�xGGG�ɫ/+��`�+�VOW7��{�����\:{���N��$�=���:�x�ɇ8��w�{��X���9j,�nC�<��O�/|���yF���;z��H]����ӿ�y����Yؘ��62����o�[�ű�<��o���l�͈���/b�5�������>�Y����ܹ2��G?�w��&i|�]5�����Y��ϾBri�����^�=����jj����?����?!����o��:q���@o7u\�~���2��+K<t�
��N�
`n߼�[o�ə�giaQiYT���-ҩP�d:Óy��{���&ն��X['���[Q1r_��*ZQBK`���8|��ݝ�l��"����e�_��?�����˗[������dZ�d�����A��W;��E4�j�zb�n(d��7��ƍk�B[8-&��$.�Q	3�㻤�P�ҲyL-6�^��E8AqL��`"U��j�M@�6�P���S���'��cv��k��ۻ�ʀ��3�����O���6�K��ų�cYt%e�462���SLR�D(%C�L��J�����>��|Z����::�Z��}
H$P��V�L	(�FU恵���0��Z����k�z�}6WVU�%5p�|DY�/"����L��LkC@e���t<Ehe���E<z=u��6,z#�d�P2A\�Ϩ��릭%@�8�R�R.�f"�r6���G�Ã9����*��\Ͳ�Q��lKC����ɬ�d�����&�c��U��F�hR�+�ь�������-���͎�`V���rŞPS����Է6c�z�˥"�յu�� �����Ү2^9��l`��^��O9��{�`�})mlm-�*�[�X'��R�$9~h�I��e���geq��z���Y4��� .m�:����.\��2���e� ��T��j��S�P���4K��%Wq4�t�q7;p��К-\�3��r�SW�)��pt����inÂ������05��#Ѝ�ӌ�`��^��\=������Mj��V3��G~���YΟ;�p�RZ�ik�oh����a��^�zCݣ�6�Se�RC�l���S|��_�.��j�5����������������	����\��k�����?��SS\|�=LI�WG	�X4j�����}�ܺ}��GF8w�6���:�R��~��\>�>3�SX�v�f�y����k�{l?go\���ym?>5�sp?����G��$��.������c���kċ�Mףזx��r�g�������s�m:j�؅q3Y��'?�˯��Zh�G�|�wϼ�� X���Q�������T�X:�ɇ�b�U��fgme���g>����yńH�V޴0w:-���?�ɓ'1�̊ڗn��e���S�͎�fU��f8��tES[[�G?�b�Dx�n��=���_��}���s.����RD�	jk��D}2�/�N311��.^�([d�NX\����
�^�p�|2��b�9��j0�t�U��Z-�9Ra��.��L(*H�'�=���l^	V�>'n�	�Q�(g��n��,��-Ej��Եy�zdKY2�ˑ,�f���-��ɛ���~J+�����r[)��,N_;:����b4�E1�Bfc]6N�a�g�b�iJ�QK<�$�Kc��=���f,N;�WQ�Rk�v횢=z�$�--
�E`��'�v�*����*k�=Jؓ��Uf���B��@C�K��JSЃY�~�(8amv��w�����&�y�~?K[���Y6�i%����h�u��Ǖ�rx�[!�=k�{��]�O�ci.��R��Z45�d�Nt���i��-DX��"�����liDc�`�;�d�֧ak���5^�M��475��31y���@2����#�67bv��hnW����;�w��a����'���gg�T���oW�q{[������z��Z��� �\���t��RΧ84����/���F1�"����% �NÇ����٫J��+�����l�b7�����KgY�Z&e�Qt�ih��d��觡��W�8Mh��Zd��a�i�����|�~�4���,Ĉ%�4w����O��lr��?�˫c��yt�8-u5���>���޺�k/����P����`��^\^G���������L�)����𫌷��K��>��������M�Y����g�ڗ��p� ��5�;���q�r�x��J���-\Y#��%�%���>���m�ߺBS[�3c*�u��h4v�w����|x�H1IJ�$���`��7�u1������x���}�	k�lzz�{s�ɛL�,����0�jT��t�#�8F�� �8Ů�zUJ� ^2ڙ�IB�M���J�>p �߃�i!�
E�u�6�x\�C'Q��yU��V�_|���~��J �/
#��]������1%`�[��(��z�R>#���5�N�
����|Wã�>�$	����;�������/z�z�����{�FB�8�t��`�R�J =x" ���R��IW�+}�҃f.��s_e~~�s�^Zb'    IDAT�cu~���z��pXL*�~E�����
�$>���S&��!s�-�:�)0�hh���0a-�T f��u�P��ÍɝG��,3Y~vw���	�>��Z
zZ��|����"�(����^�:b{�1��X"�>�6�F��B�݌Il��I��')�QO��Z;Z1:-�����@C�W��؉�x}>U�[ 4@˿7o�_���NM�q��g3�ͨuFc ��`��h���^��k7t��m,�Y�_d��4��FK�d��d�粳^cfs�0y��M�h�b5���B+���l��e��l�l����L���"���d���%ow���U�dd5���:��Vg+Z[Zs �ťXB��B��n�����H.������ȍ�W�55��G[OV���j�m��L�L�����#��u��J�߯2��Q>����w���s��Y>șS(ejo��Ez�8yb?+<��#�y��^��Kcd��]�kj�r�ɦ�|�>���������xT���䧯���@��!�z�e�Vp5{��L��O��@K��]�������5���L���'I;�Ե��h?����ؚS.8�S�<D^����B���G�����'h!���ӯ�_����ַ��׉Q��Z#���;�������^�)��`���V��.����f^�rIѤ��_��TZ����|�ُb0����ߠ���B*��n�\�z�	����W$��i����hsY���[�dj~��O4#X���2a5�k�M�Y��1YE4��_��FO��Hɔg)bz�̝93�1|��Ɂ����𳾸���&�M3锇���������e�PX�"3Ozsb���z\&���%؊�S�k�mm�o��.;���M4�֝�lE�N<���/���t<�+���O^~I9O�\��0j�;W2��w�w9��LLNO�TW��"��6���b�Q�aJ�*ӏ�v���W����奱C���� ����=�w��Ů���ͭ0�\�@M�jё��пҷ�����1>��Ѣ6��t�a�"�x�,.�3q�&w����Bc0��nQ�j��SJ歕5³K�6�x1Qg�᧌�n"�ϳ��ʒ�ii��g7�1�qX��5%��L'�(�4�;���̸kumz�<޺��D̈�kx����,b�"�����B9��V��f2� Z�}f]|md���4�N.}��C.5�Pܼ��N����>ں۱�lX]��UܺuKedG����N�չ��_���q�զ����m����R��j\Vv��R��6p�LR9V&g	M-�K�iq�ir����1H�2���)d0��t46�X�������f~k�5B��t4�lub�iH�r,,f�Z�w'���4�%R֣��ɤ�,Oo�0�Br-���Ec�A�)M9�eӤF�e�H�ݥ����]�j�hM �"o���:���{��r*�M2���f��zWZ:�{����Z�wn�dzz�����V�?O�)�4��?�#���o���٧�d��z�8~h[�K|��>�ų�|�2�u�\z�mڭ6�$�HDU�/���Z�����4=]�kl����؃\}�uƖg���ù������k�����+o�Q�;�^��+34�<H�������Gy�?"��&�231���l
r��1Zj�����&���}��������#*���w��֢�.T�I����;�>�N��s���)�`x�,V�PI\�U��}��jV::�����x���ܘ4%���Ec��]K�߭4w�\!�C�������3`.��{�D���,/`�א*f���&h�P�� ���1���\*��F�7��ހ˓��ұ�0���Ɯ�+�t���փ����&�c���u�?�u��)9И8�Z����ר+'�$6h����W%�f#�b���9�n��:�V��ۮhwa�n��a#�����ر*�jUp���7���?��2���	(a�d�ʀC�W �G�G�u�+�V"�T��V]��j�"⓲���\p����ch`P��s3��G���w3�e��������{��Ŏ�]#�pT��)e%�IT�⪲������+��R���-�\�7^{�۷o��������nk�>��e5`��	�HGV7�ϭ�Y٢��d��M,�U�%�J��d#�!�-1����:�B�ER�,�ufS�]%�{}�w����X�f�B	&�2�?c,���=�.�BZgGc���]��1�Dq�������x�M��Ő��zsj������F��v�B�x&�v;b�����A�F��"m*�CN���#���Sk)��Lƹ~�*/���?8C0১���ׯ*AQ:�C|�[��(�<px�C���{���&�f��$�!��ɣ��[��Ե�z�,�,0�<��iS£���0�7��xT�t%�ND�֠��c��uY�oIg���0�qq�L�����?A�ldfeS��q�~$��l��#����u�Z'�p��ӯSc�c�Eh	��jlbue���5���_�h�c0h��V�zbj��(�E���	��VI�S>|��]�N�X�U���o~_}ܵ���)��_���������>�͋g�mo��[2�(O=�$wo���{�8�=���{���6���́G����+��96z���N�V����!&F�sky���C����v`q�48�45p��]�V4�]+��x��c�ݵ���t4�p��u�I�lF�x}�A���6���Ϋ�!V����b���Rb���z��{���4���#GG0[��l�z�x��W���xd�AZ[۱Y+t�{ff�x�ͷx��7�E�*c������h�s��u�v��#�w�T��b.S�s��٫�	�����qq�58�E�~�d���E�7y����>3��&A��T1���"s��&7���8jJ�-�8�f�bi�N'����Nʋf�!�f/e)����V���2M~K����n9�jT�D�i�ۘ%>q��r�]��Mu�W�UyH�5����2�������z�1�,ح&6�b���eu]��F�;�t5�:�$�1�|�M^~�E}��k��3같%	�(]ǧ?�i���'Jj�J+e�ta(zߪ��P�RC�yE�|aٷ�ө�V&��'��s�����C�\�r���g�F(L8S��*�U㳴��1����e�f� ��1G�%(2~��.�#��r��Yz;�i�1�����ZL�i2�8��-RK[��x��qF/]@擄cQV�a��iU�z���bq�"���̆��I�Q�h�n�wo��:F����0�+I�ͥ�M[�\��J"KAk'+�4�Nb!Jj%C��I��26��&M���K8!t�%?���� ��}��L,�"	c��T3���?��O?���g����bU !Ѱ�C=vBe���ϥ����[������OߠW�����/}I)��f(����Ml��Q~�7?���<�=�}��w��ǳ$W��3�FWm=�?ű#�z�-f槩ijR��>�.�����mW��x��i
�"K��C���"�)�)�vm��KinG���f��_#����L*Y��7�RJ�)��d����p��m����V�s���ե ��!�����t"��'UC����/�pڔH������!t-=�M��	F���Z��ڣ��P͒)�9}J�|�������௭�����O��wy�ͷy�#Op��)F����$�Mp���N��>�����+�m���Ţ�P��F�����K��w039Ξ�]��Ft�"�F/3K\_���� ��3x�G�LM���A���eFǓ\_,p3bĿ�Iw������]`el���,��Wp���#��4��rs�0�V�k��h%e�r���e+��T��������X�8�v���
x����OSSM��K�W�����R5K_������j-��L��N�[	�;�Ge��|�:�S������ޚÚ(2\׊Mt��5n�-66��Lz�:��
8�	̦"�R���*����F��ԡw�0��1;�l$�\��re�Ϊ���㌧
��.5�+�3g��"��]�bl:6f�*7����[bo�����^���j�f7�NGY^���sq�G�����j6�r;�e���V�6h��T}�R��W��L"�믿��fa
������E,v����Z��FFT+��ȋfC�WG�Ŭ|�vg�k��A i�:�9��` /����ɑ}{�4͎	�Z�[������~�j}SӞh4N4�dffFeR2�+T�xHˏ�GU#��j�2eH6��f���s��֘�}���v\���{�_�x��|�o��&�Ë������a�9�(��{��6���Vװx��E���C�a�N��F�J�Y���f�X�b�ޑ���i
��E]�r7�g<R��ӟ������/c��3=��̝r�����|��������oP�(��Mݤ�RV ��~����÷��uj�~�^�N"�"P�l5p�c|�ӟ�埼FkG;�+k�)�E�l>�ꅮ��N��[�op��Y>��{���3�������+_�*��<��Č��ч���ϟ��w��ُ>������^����xs�{�nnfi~�c��$��ƙ3��54ą��9y�tVz���g�`��7x�����/10\KCw�fl� �����M]#o�X�ݹ��_}v��7_~��FC���J��O�&7n�������7���:�lN��T[C*g߾������V@���[��0zQ{�����!����~z���,���^���-�_�\}m6��Z���O*������3O>���4�A{�To���BW(qὋu6����P_��2�p�{و�Y\�$�ɫ��ޮF�.Qgq׸X�opgm��.���B�@-�Z���Y��V�s�6��wR�{$骣hvc7��lf�u��sI��
�:�6^S�������o�����q�O��@�fֲ����ֲ݆�v��b4���R%���M�'��}y��aU�ڝ*㕬mmy��~�"���7��D�!�&��Q�S�H�����GpX5��E�f=V���w�]*���~�K+��6�q���-�������}C�[X�l�2�l��D�+[����P3��nG�C�j����$�f��0|��X�dQ��l!�b����2��^j:�ҭe0�1S�_'5}[x�#�n�ҩw0i����ɤ��-Oh��ēc�z(���A��iW�O)-�,3��C��(�J�i���o��/��CU9p`�/|�����bV�����*��+T���q��'Է�J2��]z���o�~j|�\J\���4�gϐ o�W�>��{�ƭ[��M��pLm���Y%��XS42�S|��=���5�� ��!����"�wX�����K�ߋŬ���<�ѧy�{���k�v��׿���>�8q��qzF�p��Y�g�pjXmq��0���ؼr����en.L�0����(C���u|���i�n'��n�l��ur~r�O~GKHcGw��3q{g����{�>��G��g�ǩ	��e���<2�����<��Q:��8����g�?��O	��������g��ݬnn�?4���&�.]"��� e��C���V������Q�~p���i���Pu�`P�b���!��������ԳOs���飫���ȯ}�\9u�7�
CM]���+�k��m���:N<���i��y��G��O^偣G��A٩����7�r��\-nb�10܀�΂�g��	p��m�bz�K���am��br������dm.B���ٙ�棄S(��}��z�ish)�M��\���Q��6��=�������W�__K��z�A��lf&gfT� �{��Qzz����Zׯ]Qt�_��_)@1h�*1Z�j�d�=��1�I!��r���ƹkh#)�s�4P/���<v��p2��ܚ���ɱo�.��F[�6�1ƶ�i�ؚmt���+�s�(a%����u�/��.�b�?J��L��¦�_�s����G&G%}#���L|�6,��^fw���AG1��n1�X��Z#�RO�� =�}h�E�.F�A���N(U�(z�`�(�@������c��;=9Nx+���5�J9�����'��rQ�֊�p�Ƅ*����ǈLN���#`�4c��D�f�:��;2H:��6��M��R��x���'��>�D83�ú��i`=V��d��sN��L�f2Q U,c5Y�.��:�Jj�D�O�	�Mn�39�]��򋷱��8�^�pK�.�UT��禐������������}h�:e�"%�T�j^X^bp�������ŧ4
��;o��O~�����ad}�f�*�<��kj(�*5]�⧻?�Z��R��d���K��ϫ�!����AS,J�4;4�'������+��\�������Uv615SqXI%T=�n2S��gM%������څYE��r�۷�1?9��i��Ə^WR���|�;�nq�g�8�6�K��<}�&vwu��n���>«k,���������릥%@<�D�]�Q�N�2��A^y�e��6�w�P����hee)̭��y7/��Mϑ���l�a®�\�6�����]���jkGp��Y��88���ȩ}��~�1��������2�k�������7���3<x��/�a��A�j"�{G����̙�j�B��2�hmoS��x<�]Z\�?���P[�Z�dx�o��o`���ۿ�K~�ӟ��^��h��B1��#�٘_��O���~^}�[�ml�k0)��Cȕ2���?�kW?��w��R��im���:66׸9}��_Kޚd�P3��ۂ��fll��u�L���bj�E���m#��\g}!�!�"�ar�%Q��3��l�|�����9|䨷9p[L�)�ڛ�u��w����6Z�z�[��L�ddiuU� ��ttt)��d�j_��������3ɤڃB�J�F!�S�]1ŉ��iZЖ��=KF�Lߜ <��#�gOM5-�bN��$rfVØ4�"��}�[��Ee�'�Dx��bg��]�Z�x2�MiJf�H�y��*g�,��q�~��-H�����Y�0ui��B�g&g7�R��ƈ�P��5Gz���'z;�s��a���	�C�m�c�уt����'��xQ�S�p��(��G{��0��UZ��e����+<���<�أ�� �>3��+�$M9���A>�ɧ�GVHEV���T�3wg��;s4Y�|��Cl�ck�uh�L,-BOcw'{G�ID�)���4d5fb!n�Ct��mo��$�:6������).LZ*��If2�+밚�$V7Y]%2]�6��w���<Z��x�Gg),�E�2��:7}/k�SJT��:I%#lƄIs�7<�[�W�2G��ɥҊ�_Y]�kW/{���=+m>B5�:��W^���>��k�928Ag��D�"r{�^���Ӵ k+ ,@m2���`���J����{��w�������.��V�F��~|�3�3.�n���O�����ؘ���:�+y�w�x-�f�)@"J_���r`6�X]�����v.+f�87����Gt}���I�n��\��UC�b�`���ݢ��P$ʞO�o~���V�^�b���:��w�f	��pq�2�=�.J�<um�l���>f:f�'�A�#g��Ե���&�i��p�ݻ8�ĳ&�v��-t�\z��|��/|��7բͦ������Tf{��i=�������v���T�Rf�J}7�H�����Ȉ�I`"�~��I[ǥs������5�j��nɍ��s�:��8Jlk�=�Zh��`�h�;��ci� �/��8s�=���Y�r9u�4%���&%>�f}�-�Vr�0;tj.���q{m���c�}P4�)�����]�sm��~,��I[\�zr%3�l�$ٜJc��br�'Vt �n����-t˓8�˴Y��YD�S���-�(�p�x�?����.4&6��!ul���AJ@�'����Ue��do�LN(����/+ǟ��ֽY�6�Y�,���G[J1��A�ߌ���m�(�]�e��������8�Y,�&m�\��r,KJ�;L��A_
�Ӥ0�5$5E�B�L'7�����Pzg��6F�Xb#��+�|0�f��G��O2/Q0�q,D��L^� ��Ŷ?    IDAT#�~�����_�c1��>=zOz��ޏ%�fmaM)�٤!���Y��X��'����d2��I�r��7n��ƓO=��PZ9��^���W_~��}���ڳ���O_��L
H�RʰoO���ǉl.�
��6?}I�����ǩ3����D�'ILMP�!��3��l�Kۚ��C>��U�.�g*���h�����z)�Wq:�p�Ml&����̨�k������J<e�8ImDY����x�Z�>��>�i���c��D�),�R^��k��e��H`��q�mĢ�
x�N+���Է�`qK�׬�U�w��es+DϮ>��2ӂ����$���ҏ�η���R��D2�>�'"�x*��?�y�6�B��Lc5��U�w�PT�]	�$���<_(���{�%�׳����v��jkk�����^ևxO]�r����?��U���^��N2esM�ż;��٧ư���g�(�bܸx�A��f�f�1dZUI��ė��n&)�G�q��(�Ő���������V#�tu�(U���T6tM���2Q����@�P#5�N2�-,N�[9nLŹ����Z	�zѲgM#���'71glL��P���CB+f���u2swi5Av~����RMf�1l.+�D�H2��ί���wu)�zOe�:��J��Լ�#G����U1J/�I�⌎���ď^x��ϣn�h"��A2%I��5^�"�M�ߎݪ�*���w�_#=��=Q����l&`�^�4Y]���9�ż�p��!Z&���ΐ�qc�-O�i�`h��y�{��)O�Xbe5���,�u�l��ڇI[�$Ż�`dnr�ŉ��|��$��h�-��h��8�;8�+t�4:��3Y�F�Г#������wr��h�륨+c7��2T&�&���#O?�����M����ys��v�a�gz�'af�A  @� I��I��*Y�u��e���-��d�je��%Q\�@��0	�C��}s|s��睆�� `WuM�t�������;O8�9����e��>y�s�����.ϓw�M��d%����}�+-ee���Le�k��d@�����_�4�s�
�j^��F�c����(���[/�1B��ZҶ�q���n�p����hR�z_�����c��
����?��q�[P2p�}<��	�]�W�Q���^�D4����.�������ۯ�=�?~�8pa���P�4�.��o���y^���t�����{|�����e��3r�}I�T��?��������8:�goXڻ,k;XZ�¯�k�z5��b�6���[���OPd��r��!�Z�$+{�kTQ�]�Fqzy��@O��4t��6���8��y�>�E���
>y��O	h��H�_DK-�8����=nc��.zk��_�'�#�Ԡ�>���G� Wױ4��t6��v5֎���QcZ^��K+�]Z��O3^��X��Z�x,�?��+�\&.�x�uZm�ş�����<<���0�B�ʚ�����dA�!�Y�oi�\��M#�=`�u�6F��y$���K�/��GG�å����p���9^��޾sdb��Fhu�\v!�%����p,���S6$xnEF�G�UJ�,�λ8�x
����`�A7R�1��GmkrӅ\�c1?�� B]蚈 !*D� '8�<�rр��L\�^�c�[Ƕׁ>S��bcg
P�mDB�fK��m&���<sqia&�D��jc��1��}X`z�Mxr�Vd;����q�l� �^�,t��}4�j�.��:��f�&N/-���6ͦ���zm>A&�c����t��J^ā���g�}��_�F��W�C��28���6��Oϣ����e�
LU`�3�Ox��
A�y��IUE!�aj"ډ���t$������
t͇,�<���`��m���W��i=v�9������� �|���hK9؂3S���v� :
11�*��(q��rU@>^C����!��X(aժ0��'D<Oyܮ@��x냯bv�,��EƤR��N����M4[-|������g^�t�Q���?��������gp|p� -S��4���ܹ�Ss#�w��-e%Tw֑S����>��ݧUs��w�����nc�L=j��W�(

�|��_Ck���.2�����^�Z���+�x��p�C�bT��C�Y����h���_��w��*&������'Oao��x� hsX��!�9h����	�z��}|��k�&�WW�t���-4��B�|�L��fMjr�2����ci�|�(��Pu*U[�����������}��9��O���n��`�p�>g��#���7��}d�%�`}��^�wV�;	��OCm6Q��1�i�h��0=7��Ôm�����š��j���c8m�0��6 q��zb��3��Y��������:xz{�v���W����A6L�Ȑ���`�	��>Δ3��f��A���&5���2�,V�\���"Ԍ
�TR�y7���wa{>ٟ>���Y*��N�Z�G��ٟrv�n���Q1W���o���+Ҭ�s�S� EA.[���8�T������1~R��t����G��#���r��9��_d��r������E�v�Ǧ�D�"�ڌ���`�K	�����iӑ�#q��&C.:ԛjV�sqjBh��m�)�p�l9+�P�a)?� ������a�U����C/^���!@�:P�m��z����c���f1vڀ��CPbԚ>ݰqcWŪ����+p�4��p�Q�Y�~z��NQK�������A�߃���U��#Mȓ�V`��%���g�kM�������3��AJRt�Ǐ�!W(0�wbf��!�Ь3e�?��`Qtr;9��!a�&B������I�[���P���&�ͻ!��=C��>2}�fΠ�ZP��,��&�U+�E!r�<��?���T���H�Z��V�EnyK��A*�!��T��qg��OvDנͽ�W�'�`��{���cx[,-�A=��J[0��%H����Ptjx��,��9�>�H�N*y����5!�4|�;����2�*��jZ�6v�vx���oa��l�A����&~�0����xx�>�wv�!+\����,N������ 0'�(�&V�b��S+9|��w�����F�{t��t�����／��[p�{(dXI��fk�Ư���+�K��ރ ƨ��[�񏏺h�.a��_��j��GVP�=hb��zO^~�~
�M�^�"���oރR�»�����n�gA�B���H
Tq����&�M��u�n��q�ӻ�o�q�b�b�+)������?2��0W$b�*��
8�0�ׯ�GA�Q�D�H�܍q�y���[,Oz&?�|��$y�
	A�N��8Dyrc�Ed�	2����Z���~[���+�(/��+kU���Z�;�l�YS��C�x	V���*$QE��£k��&g^ES�"5� �}��]X���Vp*ob��a$�pF�e,����>�cX������:�@�Vz�$X�F�VΟ���%��J �O��Ii}�!��R�K����9|��ڗ�rn��!�����\�h�)�!ॲ�'7oa|r�ef	x������o�r|<;9�R(�.�s��/5�����J���B��������%sf��jh���.�6,	J�5���l�<hb��@����S#��a�51
q�����$874�كi;��RV�A����@�k�r��Ć�w�J!����v�Bш�so]@f$ �u9	�G��� 65L��>�� *~�#J�Z������u�>@'(�2�`[rV��c��=\���v ������Nm����4^z�F�Ē��HX�2ލ�M�f��^eV��<lO��T.%��W�����m�� ����tľ��r��%��_����4Q�a|����lrs�!�����z���&1`�;��E	����Η_����w�\J2�k�C�y-]���R��/x5c㠋�;.>9�@YxکW��&�y'�n��Q����ꕯ!_��g�}ԭ�A�n�޼�Ѥ�^~ú���?a_`ihu���}�y|�7~�疱w���.��j1���n3��/��̂�Q
���o��/�;��;��_�u|�ч�X]�!ьd�f���������[H�t�ȊRZj~���Gk(D޹|9���QES����m�8Z�7>���8M�+����Z���p����9Q����j�=��,�G��u�Ѱ��GA3�ܮ��ZE�a�ċ��E��a^!�B��}�	��X�����d��,�R�0���9��֛�;��gy���j�q��}�r���k�D@�j��8����������6MC��Θ;n���sgg���)�2�!��ȓM�=�� t�9l�T#��k����s��!c�A"��5�ץi� /O�|�@vT@��!�2�!�ٸ�.�:a�"�� "Y����u<����15��!�HZ`A:ZC�S����dr��3̟���G�����8�be2|�"<|����e�Z8���vШ�y����G�7Lj��)���S�����̒�˥f^]39�% &���)W+�u�S���{�����/��/�t����0;u>���>����/�O�}�/]R�*�:����?��c#��׎��{���<@�b��Û����h($"���}�*����E���.�[��+]$�q��ܺò��1�v����R_��u4�w�EL9B��c��)�UW&q�k����	�L�J��	�?�`�����a�4c�)��juq��#�+���/}��n]K>���6��>��Ky���q��v�ƙ����g���߆�+��{kD�bp}��Ro�uã##*�G�F��wn�Ư~���?����7&	��f�`���"~��_�ݧ���Bd��~��{���o����q�9� `�ZE�sY������8��x�	�v�ie�q#�g���_A���w R|l;���N%L��҅��j��h�����o5ѭ����%lE�Z����:Oo�dU��W�`�0���m&We��>��u�G
x��cnq�{��Ds�1��.�%�{��g'�:"��m�������������;���?B�V�
9��R>B�S#x�+�ar(�^���ލ��X�� e_ĵ�\�PPD���Z��&�����B�����œF���,ξ2�Y[��p�>.��˛}�ʋ�.��va�j@U�;ؿ�o�u���\q2���.��>�g7a�w���2�C5�JB--#�kU!�	���;l0���l�IR�d'w��-���q�G&	<c�!`����Cf4���ap` 5����G��b�J&b.�_ċ� �$�(@��ύp�t�O�0�e0K��`Z���mԭ.D)���F�I�Y�(�-����z
0��$�!�<�G�;�[�-�?���C+o�q3,��EԷ�xtkQ;���W�#��<j�D}��[��\c�X����J$`��v���n��2V^8���eP%���LO�w
�._���
hN��v��x��l�:g�T:�3���F0:1�4����<�S�c1���0I�̙3�K����ﰖ6U4S�����ڣ����^unj����H���9^�O�=�S|A�3�X��bv1�@��=pp��i���$��L	x��&�+��"=ƷP�_ǻo\�����S!x}� �q#r_{�u4���=ڇ!����n�(�9X�W��6z�
�^�3_�c��ǽ:�g�q���
��ށ�	�l�x���ޞ��xSo�
�CG��DR �>�~r�Ch������p ��.dI��>�X݁v������^XFج�pkCAϷQo7�rژ^���w�@i�̦	�&%�%�����ho~�:F����+�Pzc}?�����'7��w�C�Y���"��p�����g���_�.h4�`*G�O6qxw���[/���`}"�h	d����!����K_~]@��Ô�\��8¶�Dqq/�s�t�(;pE�5��D�dO&��<�v�!bY�&���UG}����oA�WP��p�B���w�.��&��8��lV��E�.�n5Q��Ћ�z�L�ϱM��	���b���[���7?���,t��%wG��������}LMN`{{�62 �?j����i�wv��J�?�����0;.�Ma�|�ɍ(� i:6Z-u����Y�@Vva*	9A=�c��Ķ�F��/N#3@θ������V��o�X�v�%�sC3EDA��ݻ�HH�y����a�d�*Z{6��=ƫSC�m�frE���=��V{�����{��H�t#����|��-L�N�L(:$�\�A�Ѩ3)퓏?���8vv� �?�"��m�0����˧pay��rUFA��=T7vp�hSz#��QEG>NG
ے��Z��0>:���U��KT�jb������(��&r�YD�7��k���:��*��s�����ITY;<����[���e��8)��n��3X�� �:&�o�:�Pд�ȗ�X8wS�\	��*x$�B�w"9H���Lg��On�rδ����
�����_A�T����R�T��UÞ��P`Oej�����{c{6;E]<����	>�v6������?ǰ���o�ʗ%�|����>[�T;>�$Q��zt��c0a�n�vV�f6�B��U�~������8�I���;hcH4p�p����"D���N��,�ͯ����BpZ��~Gv�;�se\��+�O
��g�� ����k��p�Lc��7�T��J�0� ��͇���H�f/|�0��O�\�֫ �~
���E�fǐKĎ�������[L����/bz~A�ݓ����HE�$1F7����L
$�������=�|�n<���J���`Ʃ�Q|��1PP! ��Wַ���#��,�L����a}(�������"7<�KWΡ�� x.W:��ݩ`�&q�._� �hC�V`G=�"�ۋ�/k0u�y-1A�yX��o��^m ?u�~}��D�B�h�=x; <ù�<��2��+8T�u�����7߹���IȚ��;*׻���A;;�x���`jr�K��N���4��� ����J[`�����P5",N���++)��E�D<�[_݆�����$
��2��|���z�^��3X85��������l��X��P>���S�
6
C찏Æ������)�.C����+���{!:Gml}��p�����y
�d��WJ,���cЪ��1�rf�33+��o�ڇ�T|���Q��/Aճ̄'�O>��S������;P`L���[��Ec�#�U�x���kT!`V���42� S#sr �۾�#���K���l��*�q�UIP.e1=5$�Hĳ��1v�{��	&�'����!f)䐰�i�֓6;ԑE���F�"l��mW��ք���<De�	}Iք��W�Vv!�>ی�g^'�R�v��*I)��e�M��P�LSミz��;ۜ`���u\,��~e��V�kk���{�˧�too��;���5����-f�C��@�"��	|� V3=��Se�4
��9�(ba~��C��k��ų/�͍m�x?�+p�ɓ[�b���88�`}c�v�7�G�ae�,�g�����Z��?��!��H��f�4Y�� T�Vqyi�]�ש�ˀ���z�uC�g��4�0m&��#��*�҅^��K��#Nh��j�Q�ɘ�3o\@qZ�Yn#�-��7���j��h�s�ae��J�T2{v��>⚊����
�|U�, �UC�����=�8;3r��!r�v�˥�.����3�[�g��n%)zX[��B�$I�ÑY����������S�iӜ �/�_���s��x�(eU��I���Q����G1&pvpf���w�,a�Y�^���p+���!���c���X�7��������(f���^���?�F��_�4Z�    IDAT�?r^n��ꩊ��=��z��.
S� �g�w���,4!���E�>��6�(�b��X�����&.bx���̃��)�,G�ǨVk,9:2�YY�E �7�?��������ν7
Xh�'�S����H	��
J	9=�.��]�����������4�n���� N��ZG�����9,.�C'yȌ�0��-l��X�41����I�f�]��Z�Ǉw�����  '@ؿM]@�(A�r�ժ��~g�F���D$��S�!�������`��V��& �}T���{���Fs���^������)@�13��
ԍ70�x�����B��*-��;ܧ䞸N*j=�$�O�KLf[�����0�&P�h숕!񜾃��m46�����\��m���\4�X�I�2[����r�Y�4�pZ�
2#d�L�fI�'h�:�p����C,N@�/��s��_�G�Ё���0$��P�`�D6:�w��k��yE�.�2��I0�&���-q2��Le`:�Xן>�,��d*�	��6�99��s��>����@Q����q��U���!�kΞK�rf��ǹ��5UG�DHF��G���340 CS����������W&''�?ǰ����'7��UQ�qxT����5������=�3�x����6(R��꼁	ӈ�@�Ce=�=8�C��"rj�{u$�*Z;U�vj��"V��tz(2B/�pԮ�@F��/BWbd��"D��N�ZUc:�^<����������d�=�F�.��0�4�3��z�����K�����)2�*�]x[1t�ӳ[���@�N���h�}�.L��s��H�mE�砨xwk~�ʕ+���a���i-I�������{��<�O�&: U�kU�Oy����(��سx޵����1��qa�4�z���*T�>g�4+{��%X��QYAh���j���Rg���V���4�=<�@�y��,��(�H>1��Ml>ރ�������E�l�sЅro���0���0VF>a�u� ��u�6�aP���W�Ʌ�>�LO�p���#t�=|���8� ���󱷳���������dH�̎e#N^]P�kx���,�H�^$gֽg;��� c��02��� G�j?����z��a�OMa����C�v�`��Į���J3�G!�}d�}G�Oo���~e�2���"|��>��t���W[��_A$!�� H*�a/ck�S�
^����0�<"��344�W�P�ᥗ_Dix��*�Q��\6�������TC��)�$���o��o�у��Ҡ���rq�K�RBA�����ɱA��J�,�f� c��S�*u��.�3yS9��JM�Vv�A�怐h�S���Ԏ�uxB �lB� ��,�"��i�#7�b�����CPG����P%[��Щ9P�e�� ��,�W��7�Я#��Q��160��J�,P�w�I�AL��M[: �^��n��Vr�/w�e�+Ut�ΟZ`����|�Ѹ�5	�4�*&��"��2�d+���X6TU�@�"6!V.�E�x�$j���ryt�����߸8I
#��/<����'7��򋒢���f�6�o�2�(�%��˗.��n0��>8�,�T[�0�S�2r:P#��L$V��<J t���5azΎN� 6��B��$qQ�ڨ�����K+�d$�Q��b�[óV60{�4���Ī�V���>n�G��!�^EP��o���S�bgm��5M�g��HC�W��F�f�} �J~/���[=��� f��9z���f7Ϝ����Q,}�D�"�=��c�t���f���Z}.=Q����|��13=�����u��)N�)855�ׯ]d�#��G!�Aek;���,�8��丆A��`VG7�� u�fZ1��_�
9q`��4�n����6F΍a��,Ԃ�l�N�O�ww,�ܓ�L]�S���!v��$���-<����vó/A5��rR�C�*�}��C�@.�PT��{hvk�.����Ayp ��A&�A��xأ�u�Ɨ�x�����J�l�o����#�����'&���cz1�
��'S+���x�+o +��	�J"�pc��}J����" �l�!�+6�\�¹�S0� 	��1z���vG�_(c�� 2�fـ������� ����KC<ǫ��ӛ�h�XF"�e�
���XՇ�@ja"����(�8K�U����j3�{vv�rfa���UʊIkzuC��l���g,NL&�?��?�/��q6ڧ$r9�*O�cB�xv��ˢ�/ #��|����w\G^V1hf��͗�8����\�Hm"��b8A�Yc��/=o@4��pj��!%tlw��Ɉ��W~`�����k;��Xt����PP$�r��0�$�)�jǐ�ź���XP,$�4��Y)�$�>�O�U��z�\�#U��Z^14]��F����I��t=�{�a�z�_� �:aQ��J��'���ioRrB���I��d��8�!��!�V�����[+� �ړ�ӏ/<�>~��|i�eU?��x�6� �y|t���WΡT*�ɳ�,($C襺�~��7^SC&�I��jA#wCfw�I��I�<1�qa�.�A�h�]T��ξ��|N�Ih!��vyk������s;]�V�A2"Ի6֏\�\��c��^AX����e���>��+�]=D��bf���yt"�_�N��P�D�k��� �����ad��D������`lvg/,chl���"c��zR`E�p�/E�T
��zC$�w��6��]�j�od}�R�.3��ry�ӆШ\}T���ud"�a�z-�b+�XĀ��,�p��ed�zhA�h8��<3|n�秠�c��nPG��[xXQ!��F�їMPx�n����P�k���K0�����@����&Z� 4qaj�8�)�d��� ��#h��7�z�e)c�񴘈.������^B�X�As)t���)������ƭ[7091�d���]"�?�v&��x�����݆�����6����Ș�eQ�Q ��q�j��J���Ps�\���A��
�Ѭ�v�k(M�1<���3�K:�����X�a+���@*MB"�UՄ&���a��q�8 97�cd�������-D�#Hv�,��P��5�+d��}�q��̪n"S(�Br:�F�122G�L��Z@kt��M������h�����w�A&L�$�y�2F>Ś��$H�:gp?<�Lr�B�;�<|X��� ���@�*��&b� ��	d�^(���z�@����0�"�a�b:D�B��)A�U�91i�?�V1`�;7��AՆ���;�^#���3�p&R^���0�2�r�Xb�z�|i_нm�)�*�c(4����z���ƙ�%�5]af3���dI�v	�5�z�"ʼ)HLB$$��M��8�yO>���^y�+�S���e�xW��syp���q���ԛ>� D���@��F�P���vvwy��qRf3����t{P�WWfqf2%��8BN�;!�z��#�V��ӋP�3���"Nt�.��mHyg/���WaH|��꾅�v�)a��$�V�!g:��"��.vkn�9��0�_@TGd�'
7��V�[���:�P\�-��ux�M��#�nSY�9r��s-����G?p�-籸|�4|ڧ�F	x�kޙ�Y�����X�U����Kܺq���(2�Z��,AL�����S�X���P�\�b̲~�jO���1.�G-�;�-xb�vr�����gQ���~��p��F��W9�<���Q���DM�Q�íg�5H#KЧЃ�DR�!�n���hw�0w�>� 2���%�Hz8^�R����OA#D�6��AP�Ԡ�t�)&YÓV�#���(L�N1�# ɰ�u�j�ɟ<zLIrf�@"�� ��L���j�!��h��Y�ʹ
&vW7�87D!�`P6$ ���B	M�B���0T��!3�K-dy��B�،�D��q�<�x􌴨5��h ɐ7���q^͡�_E�H��ؾ�d���fsh�C�X|�w�H��a�-,rP�}rJ�l�(�\d�$� �7(ۥ5���I��~F-"�"�9c�$H��T.h�Z!
d�8#РroB��T���v��G�Ţ VUDV��T�%��&���м����(��IN��	)L�x���ĄJ��$2M�+�B�B"3.g�q��Xć�*E�X79�l6�HiF��`Z���J�������Ĥ*|t��u�SDbL+)y��� ��K�T��KӒ����}0߿�������>�?���8"`A�*B*�g؃��ktp��\�t��~���x��������b��=^e�HȠ�����*�E`蠣����*0d)H��1��+�T���U�za�B�=��6� A�D���5{6r�a�O��L]iVa"Y�h�8a	��p�K7�A��j�#�eg_Z���A�p�k{m�U<9���P�_Fd��gk�]��`�
!̡�613w�T@�,��;܂ҫ��{������D>G�!�q�%f҇^�x��,t#�ϳ.2�'���a�W���aȏ����ǟ����<�A�<b8٥Ѫc�����,��H�Ȯ1��Rڇ�vaU�H���,��p|�ĲX�/?:�#��&�Ǡ�!�k�۬CPu����ȁ1^���8�,�-�ŵ�U[�rsnrBi�p��C�t8vۅ*� 
#�c�N��o0�@{P�����hC��0�<�0(�����7�0����
���GɌpI��  �y���/R�26>¬z� �0
N!F�U�* ����I�@tx]J�:����M�fdK�:}��A׶���]8������Eח�P
*�āj �S��zz^�fۇ�H���"�SQ�da(���w$���������@y�r{�"�����C��%��e���2QRX�L�\�X<C�1����y��?�`�2-���
}��p&1p�2A����(d�%��EO�,�$�tYa�X!��C{7�kx��м:�J*)��'�4���'��v��������<K�O��`R�K� ���I�p6�z��8ۥ�	
R�F�2�7ҿ��ʨtL`ȕ���H�^��x�����t��ؓk����PE�0y6��G�Xd���%�N����2p���#r�4�&u+b����D!**��0�����}���,Ħ�||�3�{�������7J�"*�=y�J��%���B?���e�F�ŤITF>�y�����8](a��N"�V0�� E|+�ӱ�=w30?<�U�B�VI�.eQ�^"�v(ʪmݒ�s3a�B5��� gM%v���b�8�F=BG���Afpn$�x�	�mX��*�!��ϡO��؇D�K�*�����s�,�Gdr@"�T�5rY��;�t�:��O��؎�e���+����lۅg[X}����ghU�|(��EjM=����y� �z(:FK�$��-vy�Id������F1�j"�؉"F�gѧ[S���A�p�=G�br>�ey���96Hp�uj��1�n�a�@.��SMt<"�P�������D��+��#f@�L�䠋nʰ��P�;���|h`zn�.Ï���d�4��f����7"�PA??�+�>i>|� ���}/���gA�ɱQ���~��3梬`ll
��a]ݬ� ����4�L��A�5�$�!&���f�GR��`dr\1�  ����b�ު�@����	
�l�Bu��
*��t��m Q �YD4����&����BF�3��'Hs�	�e>�I�z�iV�8����+��f�R�IkI�6K��>W�h����Y�ր9-��!����$"�Q��#pC렳 �,�|��E���/�}p1���R���޴�_��A|�[�����:x��_d�г����M�2�T�'$�S��uHN@>�����OT�(���!栆\�U���		?�M�����9.�D?�֏֗^�&�-&�4Q�l�>��KߔU�ѳ9�\�����ޞ����rO¬/«��y��?�Aqh�[�B	G�v��Ղ,�%�dm��H�d�N�3:��H�Y��N��d� �݃��M���Y�zFrB�	~�C��eS��XB��t=�7��+�kAQL�P�j|�T�M4}�"�F3(�)(��"A�bu���v�f ��Q��EAE�ւ�w�x
��\Bi�J�#v��B�Ն�nb �A)�a�!�䲬`E��<��˥��'H��A��c����4FF��*�	 �K�v��tߪ5Ғ�f�o[�"g�O#k���]�q��i@cXVjTBj<�`%z�3 Q���TQ���8<E�E�'���`B��2�B�$"$�tF�(8|��{H|n����\>%޾c�����d�@�*�,�p,RL
8k�e4L����N�Sy�v�������<�� �l�G,pbJ�~�C�,��t>�耢�
j|v'i	�֊��t�y��j����.YTF�AK�㙉Q�n��02�DI��ʔU����Z�/�|���1�6�O�I�R�����˔䡪�:�v	���D���l�aÐl�Ȥ(�[��`�sn�x��Ǳ��f����$�(`Mt��Rʺu��˛ĸ��bPy��~��Q0��(i�R�#��I�����!�<�BNX��){�}L}Lz��{4B(1�'���8.3s"
��Q:��<���3H�U�K�8MX��ց�)ʹ�1��I	y�>�Z�t��_�)��9C�I"e��'*�t��i��{�gK�?����Y%��@� 	�?��!�=��7E�t�릵�~:�����v�y���5�U5(i/QO�YJ_1>3�B�۲���~������>�������Կ��D��gХh[S#m2k���x��B�3�~�!IA���ZL��$�t��;����j�P��˖�k��[>fǧ���߃�hn�`�T��� ?g�!�q�H�jdsߎ2�e"D� �?1�YT!!
CY$2E��z��'¡)�l�n@1��QV82��,���tݐ�
!�}�3�9����������J�d�G͎f�9���C�G��*���Ф��^��Id�}f�T��IT�b��%M�AB��Ƴ(3q,> ،��0�J�?�~�
9�A�fn"�mSO��J�>k�BґhxD�#$�Y�!s��5��Hz���r�zi�����T�spE:�"L>eX
+�U����DvB�|�(|�;�Y:pR�TvԦ��x&\����IY	���9���u��D�#�(�s��0�{��p���4)�	�aB�?�Rr/ �*0��3��@}�Hd��,�Yfz��,���L.���vҽAٴ")�j%�^��,oȏ��&N88���k"��PDQ΢z}2��˓��z�a��hs!�ynPB- ��I��hN|cy�P��xn��&ϋ?/�Ҟ�D��BJ��\� Ŭ�N� ��)�� "�H&J�yʎjg�qVJ w�)�P5,��N^G
���K�����=��@��u�!���K��Ǥ�q�^����S�9Nx�Vfॠ�{�ϳ�P>�֘�)z?W:2D�J�4�!�2�Aj�:���Xj���8��齤s�A����O&K�����~9\8���++g~����������0>5�k��gay�m�iC�A�}�N�Գ�<��q�/"�8H\�,&�1�z�"r�hﳉ�CC�,c�<đou� �f��c����D��Y�)�4!D�1��	"�@DQ8H��،~�p谊���bR�	w��|�qyt��|�@싐c���*��*����11��E�ѥ����zF�K��nhUKg%�(���B,[��� �2I�#|S:.t�z�X��G�ЋE
b��1P�*�R�}0�x��$`/�(��:�(^�m�E�Pț�>��J�$��s�K�T��h"    IDAT�J��/NY�Y�ݥ��0�Đ���!�L�\�0D(�	A�����s�����D�:�t�$`�g@�d*NNX�,K$Ҝ#�8� ����i���'5$:�t�ϫҚ�r=���0�ўdc���D�D�s�Y���ɕ���0�)�����'"�YR��d���_�7)��{�Գ�D�/da�|MtEJ3�n����]����tĄO%x
�/N}ZQS���^G^�O.�g��'`��aa�ĉ�0UU����-#�ƃ��S�J��'D@���@�K���F���TJ�^*���P�%&H����Jp@��KA(�7��/��O��t����r4m70��k���Ā$�d�'���=
J�e=L�f�O���>e��3�$%���(4�J��2��`�΀�k� ��.����Ot��tJ|p:�4h���ꂦrO��݅Ӌ�:=���k�~�����@N��|�^���k��������������QJ�7HJz�H}��UV��#^�<t R(ț)��*&�Y�&��>|�CS�C�L���G=-�零jdeGt~Ea��S&��q MX��YG���@8$�%@lE�V#._jzq"�Am)DL�E�D%6�S:���C/"0����1%i\���#*eh��8j�CB�k"�PT�g��3�%P_���%�&2eU<�~O%}*KR����Ⓘ���s�>:��@Hx9;�RrL�C	*S/�rev"�����P��G�{c�����,V!q�$dl�������\�INUz�t�qFI�ZR�Q��~)��Ϙƾ�AM`�����=�����i[!��;��V5)�����P #�{���;�������#B�6�=��J�K	l�#%� ��"x� Iͤ����PEdI���в,d�E�{�3z�5���iI���~G)�Q������f�H�umD1�[�J���,���io��#Ylf2:kr���4]��r6���p_5ˡ��������s�3`� <����@@�c.��>���i�=�E�L��3��`H�to�����ZZ�*h� s�M��}Č��	���!ÀG}��Y,!E�~�#"Y���Q�����.�=�s{��f�_U�$V~K�9�p��x��I˛�tM��`����̜~.�{|��>/-Se�A��E��sH�����{�����&^	eҤt�Q�M��a:�-
,9�x
�f������s_4���G7n|'��gN��ns��"6*'��Û��f�f����)�2!�IW���."�Vb�xr�&gT4�O=3PIN��i솲O"�(�F�LY'������ȃ��<�J�qdF���	Ӳ���TZ�4��\N����dZM�HrV�B��F�����,"�OY���d&$�2��B�$��uB�ᒺ��`@�s �9%����( �/p�9#�9s�,G��1��	W
 d)E�E��T�׶�Y�L�BY�%��7U�yE��D�.����"�~R�UTM���	�(5�<_[@�f�Q�/��;�Ϊ�_���͙�I!����{��H�7B��!�@0�� 	%)�E��^�%tI=@z�>sz����{���q�&��ϐ�3�m��yֳ�z�q�EKd0�T��|�t�Kp%�!�����;x�H�b@&��d������K�QU\�CoOrE�x9��(#+r�A�N�ޒ�J�#C�h���
u�b�R�h�iȩ9�
�~�"u������p	TM�3[B��I�8�[�M���?�T-d(�1�� �2�}IaB"8���"_ �F&9b�����%���&�NiL&��i�(���3�$%e�\�`�RI�T���Y�l*ߪתP��@c�4G���%׵��4M�2;��=��0�` ��:�}fB9�u��sY��4���aV���ZRUm�`�VsiE``	Wl�ȫ�t�GB�m�Hf�����YA�ӚGG�k���I'C@&0���;x�<[Z�E��7�1�g�ϲձ�/L"C��{��Lp$���z�3�q,����T�L��h�7�!b�{2� �A�K%4&h�y���qφ���]��6��h[	�F~��t�>!%
�M�Y1ާ~�,����Dch4D�׊e_#��/XEkK��A�Ғ�3�ܠދU!'j��$����#S0�?n�4� ���B��d $���*���|�&�"��v�d���a��.\���@㌢�wJ�'�1u���Y!�X��+�r�W���nb4�'T�k� ʏ"��=QG0	y"dy�7P^2�1�T������ֻͬ��!�7}&�a$��Ӊ0
V�y4��Q-VU	GC�ׅ�*��iT	N�/6`,2am�E��d�-��=;_��b)kz�d�Ԝ��
J��r�50�X�W���'��J���VRT̪B` �q@��bJ�x�Y��X���f�D�%ț��׎�arA-4�/$�tv���d�o4d0o��<I��)1��u�!�˸�7žl�6_'�"a��
��Iٔ�5���5�v�uڤy}x|E�	P�(>ݣ�_��y������݅|6�vG���[$lE�	�? ���AG*;V����ua«@��$ј����*�w^7^禤&H;��t�4Ԥ"��1�<
�>v6���ZL�����6q=()bZ�����������$7�ZV�l � �i7���0z^&:���|jq�	�V˂�e���j�Zh�2��5s��i�Ov"�!���)��A3^�N�[C ��E�l�6�'�ǥ
AA;Ī��������Lq���Ʀ�PD*j����a6f_��!�����z���W���Ͻ��]���Y;���$����Ny�!q����bh�5��L�����'��'H�N�IРC��0V�U��emn�ME��4ԦC/S���6#�}B�V���a3^-�~"�̈́��ra���Hd�|�� �����M}k}�:*Ѝ�7f��p��/�.Ѡ�SC��9U��sH��P�����ʓh����ؾ�p}2���{������>���s�����D�P��nH�k�؟��U��n��/�)�U�i$R4�I�B�~æe����X���D ����8v����"JU�SY]��K�8�^���J��/�75n��
�jEw�!.uwtJ����W
L�C��
+�`R�ߥSyxш�K���}�YR�ѦZB7~{^���TȐ%,L�n��皠Z��ߗ�Q"��la�v�Ȥ ���χwֶU=Q&�6�������I���W;��l����-l��`��@�2��ϏP&5�٠S�*(��!ۛD�XP��=��[T\ߵvm�H�ɰ�y�L����	���U�Aғ�W��f��c��b>@u]dIj�L5=f��}K�k����h������_��Y�\[�-�'��|���"ׅ�GP����FISч�����ݙ|���-7n<�}��!�Gn�ˎϭg1�l���I�{�o��ք'��Ӈ#G��63N�Td�2(0w#�(m�R��)S����S�a�
�H�ƾG����O�r��*�g�dX�6�Ո�]P�we���6��⅕��{(	1��ڍGB���qS��<�Z�����H���P]T�E��1�����Kh�5�F����>�b�8��c�Z����1���Nf3�T���d�fϔ�.IG$��!^LgU��~�d z,j���D8�����T�OBY!���2��h�9�Px��z;��t�n�DĞ+Y��
��a꘷nS�쒎��k�T�tw����Sϛ��j6T���ߪHأ/��������U���i�=ڐeb{����6,�]����׀ �*��1�Q��k��3(��g�R%ct3
�e`*Gw}�|�Te3[<��m�Yز�]�り{n�~�?�z����l	��|�?"#��+��R.�iF�,� fOME�֚���D�V�jcXґ n�0���W�)�ګ���+�>WZ���X����3{��rAޭ�u�ݿ~v��o9W��f2IF�xB�{��Ň����فX4���'�I#�u&�U���lJ�Y���!4�<�1
�#G>ײ��&M��=��F���� 7�zǋ�dr�v��==�j����3��Y��LÅ_"�dٔ��3U^0l|RIt�����j��Cc�^�JWy���u�����$n����D< aТe��.&ʈy�ˑ�;��^PI������:�ڟ�*�6 ��t��Lū
@%Y	4�7�Tƪ��X������nL�^�m-ѣv#1/!H��d�ht �:�7N2
�X�h��98BV��l?�靿�&ߔ�&x�Z��j�v.wpS�8�T���K9�f��c���x�{�=Lw�|O�\��j�������$�rF|���5pp��o�/�p�0��EMf��uP���"ù g�=UXҫ��aٷ�:��{��Fz�Y�ٿg�oPˈK��J���j��l�������E\�Q�~��v\�4����\�͵��(e2rM#�k�*���V�շ_�G���%����g]���"�g�V0�����x���1��[���&���|��m����<�׺�hƆ���sš��E��'��ؤ�V��p�W���X���B�����Ai�e��3�D��dg'ƴCgg�>�����/������������{q�W��ҠA�-��'��l�\AC�NU�,IQ%y�]��v�C�M�0����y;�dn^-zp���,�X6�ka�u�[�����֮�~ᾅ��bc�������[�!z��칶"�C��i�i��uߑ͝��zM����ա�q�zb|��t\B��<�� �.�eL�ޜ;7�YR�D�/�=?��r�f�ΊW	�O[�:��l��Xh d�2 ����i[,긍��b&�0��RЛH���\?��0?��L�,��_������;wg�v)�1xh�/�c�ڵI7H�u���]p$a��3L���#�<���5	��������%SBt���h0�t׃���&rRM��g�]���ӷ�9"���HIL�,�,����Y������s��EbB�P�]�Lx虬��2������+P�[6�	� ��d��>�N��&j.���|�n�Z�#�Y֋2����5����T�&�pS�tuyl\k|��m���Z�!vI����=�z{����`b�猺y:�B�)m�9���rP�ڣn���\Ǝ°����#�`�����c�>���� �?�߆�[se�{��':�ۏ�s�=5e�O8n�>��D�Q���/���a�"Ӊ^�f̤������LF%}�I"\D빲OzO� k��o�rj���e��p��� ��u�թs�%�&�پ/7��],�ￎ,b��?������r3A�jx�Ap�j}c�t�<�,�����p����M>T���?�Vk~�ރ}V~Q/ʅ�`��4�jb
�e�;6�󦷭��J�6��^}��i�KM���\*I�^f  ��Lm�ֆo{��|L%x����0��k���q�;5���~s�M^/�fn�|f	5>v��������xj�tm�vcw0��![���+�!���Hj��|/W�9�N�}S���`�z���u �+K1���&qЙ_c��d�s?%�	zz&����;m<�� ��"֐��,\N��Ǆ�ui{4�}�ϵطQ"]�'Ϊ�B�<M�"w�&�2�Pcߏ$L%]��#A�I�L�f� �G���a��%!���T2c�,1�mo]{�e2����3�Zْ�b��$n6q�|�����OU�~>���P�UF�ɠF�Q!t��W7�D�曽>e��o����9�w�}wԧ�}�r]C�V ����!�-WQ�G3٢�X05�$�:�.�EJ��!�i�2i��u�.S��_$W��k�����n>�V����P�5^7����̆3��Q��k7qA���c��,L��w.Xl��Y1�`�?�97:e�f3T�M���#��(]+3n���1��������m>�NE�����E\�VpdU�M��۹ޥ�����J)����_�Q�2��O�t���ݤX5��ع
B��s]��XKGӟ���L��d~o[����[ �d56�l��/	e"Wuwk�t��Y����S|/�9�ٓM�t_�[�j�\��Wa�y3LZ���*��
�� �{�dK�I��d���.٨��ML����H�R�kL�|�5���Zϖ-.ڢ�$=<Q,�,f[I�w�/�/�CexT9(i%�clSd8�0	�񉼓!��_X��Bf�&������8%��~=�ʭ�#��^V��[����K�t��<��-'A���9@�\H�X��\oRߵnrF�&�[*!�%3ҳ\��Y�\S�|�-S��*Q)�P�p����I�81�'�y�����]=}h3�qc�:�y���agCŻΝ����������l���t�R�uuKB�P� {�6�����82�G�f�o�ty*|{:;�q657k�s�f D�!��l\������O�U��2m_��j�j{��r�鳦p�����#���أrP�	�%,Ʉ���2��!QO/`b�fs� ���]e��������;��Ʉ�`�&4�|����&��9G�������d��6��l��
$�4�7T%|��3�h\�A$d�^���Ti[�����l���
j�h�17L�
��p�&���wj�UM`������!+�V��[C֣��UR&.8�Ц�Um�k�H�rmU-R1/r�KHs�8=���{92���ud�$�Bl`�^�M�Hm�K��J��k.�EPbO٠��5Űǯg���DF��~au����	d��$*;Y%R��Ϧ��#c�����!�2�������nY�� Gm�<��Ke9g�H�~���s�`�*��*�&yn͸י��d��6�Z)�P��#G*�Z�c����Xۦ`�~��7�Z��?��@��C(�G_o��Ur���>3��S�{��w}�������7�4i_��;�;��.���#�oK�l�/QN�6��U0h(���2��^WW��M�-��"K ��Z�qt޺�b��9˹u�Ƭ�9�?t�pG����s��&��M�}w:T�uH$2����5О��B�p+��54�@{>kvo���8MŽ��j��m�����d���J��6�I&��"Az{��A@�����kd�lx(���j�8C�2�4��'�1�E����Qȝs?��&����9���I��A�ڬ����@~n�U��d����>:��uF�c�k������ԃ$�2��6�qR�ٱހ�Y7�$x�Ǫ���W�D�R�������<�F'���&���Î��V�(�$L����&c�l�{ǩ\,��e%.4�䈺�r9_��w�y��y��p�bH%i:�"|���e]���5֖�7oS��j��LxX=��˄����h��DI��]AWO�!����$�?��&��m�W�R)#T���;^�`�U}Kk\��im�����lqߡ�	/e����@���I�*�b�(� ЛM#�:�l�m���'�u���k��P���;�³/������ȑ�C�=�S���͘~
�&D�ª*a������̸ٿո7T���.�I��x��q���_�h4g[Wk�n!G�9�V,�\#h�_�め��lO�6��NK�
ͩ܂w�����UPF�J���aq+��{>��<w��X/G�֓��j�����y�B�����k+�~��nM��6�E�QK���{劙�c�H3�N{��Mў�aH��:LOn@j$��Ғ�"�u��:S��~�	8n�w/[
~5f��Kx�5e�B�<.��;��w�n��Ƚ�&c�(�f;�]=h��C��/9ā�!���jY#IB�4�,� ukWY��UJ��%�RW�V�䗱M�]���W2����i��(d�_��4%G��$�M���M�(�����|Yڌd�����?Ӯʮ�ɳ�Z!<�J2&�L�Mjt���Ll���Hʨ�Sh�Gј�3�NOo��D�����\�j-�]�rA��f(��o<vF��U+V�m�%0��!�I    IDAT��P*i�/v<�|�Q�W���ʕ�5ז��j���V��ߝ�%������`���$nWU�6
Y�\��<Z22���bJ(�L�p��VM2�*>����*(�5��'�o����ټ{v�x��+�?���O���R�z\SC#�.[�b���-�U9^������6o2��{A�#a�x�;�� Ñ��Ҋ���a�p�6	-���*+oq�T�a�OZ#����c��C��2 E@��g	Gv��|b����1k��,�S�sA��<��EP��f��H<����̸�j�n������h]�U+�q�L�^��n01����@���v��p*7*ycg��_����ف�r�X3k�G��]ܠ���(�Ta����=�E��Ų��E�7�h���c�:��4�'���k5��Rs��~f3�G=A��Q1p9ȕ���5^��01��ʆ����W!�� Y鬀�Z������J��1�pI���y]Hv�e�C�%Ų�r(� ���x\���Qߏ�Դfh��*��S�b�Ye5�����M�Hr�e=1{�!��P$�u�ϗP�T�J<�����f܂��6���z���>|�h�y���Gf���	w��1�`���I��I�b�]v��������t�5��oҏW���F3)-��!�/?�����9C��A\l��dLDxu��a�{���\&�!sߕ ���ikzgPz������9���`O�VP�ȆJ|�oϔW^��{��r�s!CW]�[m������f};*���ο��룿Z���-'N�ꫥ�Y�JBzBP�~r܌�<b��>A�le�A7��>͗��7w�T�Dz�r���Kx��K����>�$�3��9���g
�o�*Z�:����i�s�$�Q:� �<��T$�	MeO�!�>�`�+HPa���Ù>����b��a�~S�����t�Y�����%&Nw�dP�9��
H�<y���&Xn
�������ff�J#Y-�l�%'4�Zre�����$I�#�z{��H��a�2Y�������Š�@XKx�����E!�@���oA��� ���RX�����z^K��ަ�l���;�V�����'X��5刁��L�3����E�۷zז�k܄y)x�t�sdr9]kVI��X��4���]ύ�E��̗���bf_��P��oxŰfi�h�=î��H�N%I&d����j|m�q�L}l����9�50H����RE��R���WEK�ü��'�c��`Lk+���Ur�ph`e>���b^�0	J�v��4�0b�,+��V����Eᕗ_DK}���h(���M��XZ��(M��	��/?�/<��4R���HGl뇗bfu�f�=Md�xMW	��Z���P��O�d!>k�M���}=J��zV�`VنD`��%�����ʢ�����^ݜ���'ϻs��w}��?���+���/��2(��Dzm;�I��H3�{�q���u��rC�r���=�I<Zs�!Z�	�C�Y�_,O���;T�+)]b𐭜YTNgj�?S��NP~bݒ\E'���/r�tC�=.<�Ӷ0!�*���#��vR��L�����\��"
��|3���U䡂5}�:�ڊ�U�&�1��s_�y�1w
f���ש:����om�v��kH��q�+Fn�
h�9*v��p��B�ȠX%:6��>�V8�0"{�H�#�Vf���M�2N��������2���q�"�	7�I�j��G�5����UaH7��#����7�R������иa����KĐ)dMG�Z�=J�iq@:���&���n����d�O8����a@/�J�OU[8D�lJg�{1�!��A��P"S�(�5�p���:��lhđ�eL��m��S;_�+��u�`;g.�5����"Z�qd�)T["��|��7a�x�7aS<v�=(eS(�S"g1�eb�I�3Y��5���I��w����bْ�x��G��A"L���Xd,��"��u�1GI;�秞B#�l)2�h����l:��幺Y�J�-ܮ�ֱM�n����!|&92�=dJ�
1��������@�i��l1QGORZ�_F�����j:C-t��rщw޺��v6T��q��ӟ^kF`���6���#::��JYm��<{c��N/7��4�*+R�����-M�5^L�H\�Hl��?oԯ����'e�z2U�	\�"X�� �m��~�gT^�X�Z�Y(�P%+�\1�c�(��F�؜�ӇA�9��	>/�=��	��֒�ܦ�T,a��_d��sM
��I���|k�.��V7��럓\�)��"F�C،I��`h3eG�2�L�\�J&�bu��4P�4#9����j�N�1���ɭy�e3���GC�˶y`�n�X�����N��.�kW��������(��i���9_�{���Lk��㼚�0 �����9������L%�s���6p�S�vA�%f�
"� �c� �/!Qߠ*�h�exN������$���d�%ļ�8u�n-
Dָ� U[H2)V�\�d�ݱ{���,�}�1&n�)rq �a�K�#�Շ��݁�ja���i%�������ӹ���5搃6�!45�ɧM��eK���>�Ih���I�d�l=�X�͍�E<q�1X��k<���1��QA��B�y7�﯒b�xM��F��gfb�j���76�Q�����D x͍M�WȖ'R"�mU\��k�
[:6�V��m�Q����e���"�����؈�[||��[6�x��+���ޛ��"���]�������-[�(RȉD�#�LX�l��-(C��N!n��(K�U���?,������t,jz�
�5o-K��~oɮ�e�І�,ގU#��-�F�
G���u�%�l�c��z$���Vشs����i���#��c��Q�m��F��{�9�3<�ؚ��6>�������g
<<V�V�h��0�]6�F���?�\&A�h���p�nMEdz�ܰ9�V��p�2����9Ҏ���/�V5gaP�k�{�A�����#z&)���.1��"�@�d4.��k��57a��!JH,k�lT�����;���
v�o���C=vb�=���lK��1�"Q��~S��t�\�uq���k�R)d�z4��4��l�Um�ZA����`�KH�^qб�ǲ�s�d��r&�V>����	��'RUD �L�����R_3/�^r>F︩�ǽ���է���0����n6٣�A\.ѥ|����:M�q&��������8+V,�>�!-��G2��"���A9����d/N<�L�vw��������(����y�8�*����,��e�]��w�m�\M4�=-�D;��M]$�>�c��}���%a�K�BS�,�}�L.����}�X�ڦ�j�خ*5��U�,�D�E��������;o������w��ﾺs]*�f�;��O�!�C ���g�����	"���x+�sAM�BXMЪ"_*V�gp�D.j_�{SV_���&H������^�3X�����g9O�MW�*x
�5�.�#Tl&�0`�_ۋt�j����*��S6���-!�TYf�|�p?:�dl����(|s2����a|
f.�:�U\�U���ݦ�6b�5`�Ͽ��7��g�)ك�e���K�e?���0qr�%$��'�.-u����s�=2��ڈ����de�"S)u�5��A6����I��rUG?k�!����}�����������hh��T�����h��,�Jx���1a��5jT?뜁V�"�f�CUx]	�gJ���i�T�k�O�eNA�� *�L���ŗ�j��!҅~��b�����ڊÏ>;�+r������g���5��+הlJ�.X��u���ZK����`Pf@6S�$i#Z�����X�~���^��v� 1����-^�������Ȧ*d's���Boo���r�D���k�-���܄c�$�<�Ѓ���h�@�d��m:h���l?<�G�75a��Ëy���RI��ף��Ɏ��Q�Z#E0ka���k,���A�vX9�]�u@D��(�b�~�*��������$��L����:�a�����HBx9:�"����[v��['n��������77���}���>�y�I-VJe��c�%����t�c=�Yy��V5EP%{*�r���|E��DV}�8L5S3��L�z���.-3�D.3+5g3}kKX,�W0��{���d*����3 )�_|Oe��&�Աr�����1Ad쏕(�!�慐����	E��q�a�����Ѩ�kbR��X�d�|��u���T��)+@)hXVqm��ʵ.V�sf���U���.\S�� A�m>�z{�j�*ɻx�C��ѣ��܄L>�>Y�20��L_W
��L㥿���>����]2,�\��h�?:���d����6^g���+ U�����0x�4jQ���8Z�]'�QS��+ӎ����t]8��9<�ʴ��N=�����A3��U7�R!����Wl��6�x�8)�!�����k�Q�&���ց�eJň
������C�(�S���q�)�`��G��ِ�BO=�G|��p�T�Q๋���հޥ��I�ϣ��I��o���o�9k�A�6����H�B�\�s>2��,cu�}�9�B�p�	�d�����Y��Ň��x�Tu�Ɩ���f�B+�������8�3��dp��"�P�R�r:�f��Ke� �K�T�`���E]c��y����#��>�1��)�� �O�l"4��lz�.YeO�φ8
$:eI�#�L��b�u�vÞ��E�uϦ�Mi�E؛'�-�%��L�x_�m�⣀�%W2�fZ÷ݖ�9��I�}�1����kC��7�_�zsom�'�>z�Oh��E$�S��$k�ޭf��۔� �y���t��L��;Bj]dRʘ�o~���*@׻q� �RA37E��{�Ln<�/��!zp�p�(��Îa��=���Y��%{���Ƀ�ykݡ�#��Y �u����ve�H{U��(UCh˗q��a����b�sQDc8��6��,[�=�DH����{b�]wEeA.��濅��|���9�,�'7���c���E�ƣ�����s��>x(~r�)赓k� �����d�9l�0�k�,�B��������rU}���DX�UD��3Ͽ��;��|�ةE%��z����۠e�0����X."��C],.�*�b	���k�q�����W#ȍ��?}o��CXAǧI8��|V�0*8@��R���y��ԯ�A����u(���� �{�mjD�RB�҂HQ*�Ԟ�kA�[�F�됬����fD	Y�K�m���/1r�P445�l��T�hL���(���PHv�i���~��;m�B�!˶�p�U�p�G`��톞tRZ�b:�e_.�n5��ǐQ#0a�D�&�^Q}�E�����c�B;���=����V��94 ��_|����x� pٴ+k�â����]�>��8��8K-�'��v��+���ܻ�ڃac��%3��_"���"l��d2���g���o��N;M��yw�%s�l ��H��,�� �� ��Cw:�C�<R���;���%"1)ht�����Q;p�=�3�`L���-l&�ċA]�s��KU�i�I.�^F�x�hx�s��I�쩟=_㑭v���z2����;��C����P-�6ʏ:P�C%\���tM�쇗]�E�ĉ��e=��x�ㆿ��{㽵+?�}�I�'����>D
y�9 �Ъ����+�m咪>�yBN�_x̐X���
%$�9��n�4-�T�쿨b���m�KK��X0�ѹX�ʎi>�$�ea�t:cd5�H��9�%�%�qӹG�n�e ���r�ꞒJ�We�<�qt��h+�$����F�ӱ?Ş?�)֔H��HĂH�i�-W^�:/�~�$��g�����}�����>�@4�s{���ݽ�K/A$S0�dr�l_��|e�_�6�J��[o��D8�)]�L̐��z{~s�����q�AbĈ(����ēO<����g�:��������Fm��hX~Ȳ6�K�knĵW]�ƑCQ
��)N�P)��@2�G�r�R	M��Dģ.�T0&Q���*�G�7�/���/���"��R&�:��Pɛ�8�89~-S���d�f;�0r�0U_}��������ձ�{s�{��WQH��=��"��h��	�g���!cǀd�A�|�p~���n��ӓ���G#�����W^FC(�-'n���܈/�X��D?��p����_�@Ʉ}iՉ`�Q����f|���0���z�
�dm��a����!���ƣ��Q��on���&L@o:��׬Ė�n�)S�U��;��[n�?��1���b��C8��#��q������1c�u(��8�?F������{!���EL��&c�I[ �,���G��6�"���=�+%�~��x���q����#A+���bu�/�T.��')t��u��z�g�Đ�Fԅ|(���++W�X� �#>�	�._��/85s/�L=_^�8����T���1���]��-A�	5��/�v(�s�����Y�=&�NӬ$���`@R2�	$TqOp���)5�{��i.!͆5|H�C�� �+ ������FQ�4��>��c�<�ʋ��z��W�g1�W��I�_���ޚ�[����O�|��Sh���RAP(�Z�u�z�v����R�T�	��!�י,��!ES��O�Xf�"��ɇ���˱�	H�V�dJFJb\q����qc@Ǩ��HNMf�I $]�b�����p�N�56{L���$R�ۚ���N�c�1mp\h��e�P�M����������]�5��^��h$N;�4�Z�E#��3��z�5����:�쿟���7��ߞ|s�ގd��|��j'��c��gb�CR-�L��7�Z;�⋁DT�ߣw݋��6�!��T������,W����W_/�e3�Co�F)AT>d�E����[�Ka�ig�чB!DO>#6��s��4�9�XX�zV-Y�춻����}�w1t�P2������`��;o��v�^�C��5x�Gѱf�z��Ώ>�x3Y�L��_?�s�8O<��֬]��Æ��'c�Q#5��r��s0����-��\�b9N��/0l���O����=]���\�	n�e��gol���������o��#����셼��W_}�f܌m����6�xc���3x��Wqօa��A��S�H����H��0,�3� �ޅ�&�Lr% �2��&�v����E*է����p�5���ˮ�v;�B���_|��3g⌟M�n{L���F�����v�����Kx��g��S��9�#ڐ�Ͽ�y�ݎ_�p&n���V����^ ����A�_���0�[�_����;�Cx�2�}�Q��w`t��x�(�Ȓ F��0�d���gO~P#�9� �>7���W|�D�p^ȯ	g\��H����T�r0��ys� ӗ������B>��?{죳�[Ң��U��F�- x�n&�̵K�g��4��XL���j�;w9��,�"V�����{'�9����"^	I:__���$�)I��AǏ�W~�?⒩��ओ>�����)��x��N��֫����rY`��~���,�N�(+�}�/��le2Ԩ�1'�����1��M�/�`�.�ЕO#If*%*dj�=��W�`��?���	x4w�����h��$ey�2Z@^��o�i#��@�X���`�e����b^�K�㜱��z���� Ǿ$<28�I�^�'�����m;˻�������\��]t�q��SmƬ��#�s.6�bs��nJ^�U��c������E�ו�a�2�6ƍ�]�@,�3�>K���s�O�pɥS���5+W��;����Dt�`B>�d�h�d[����q�9��ǧM�N�TZ����c��    IDAT��|셱��zn�3�!	��-��Ie���Hӱ*���i��S=���Cp���z�_}�y�AL�f:�����_��{,&|W=?�=�f�ժ�YAR���/�G�eW_���L��YG�[m�9N�|*6�j=g7�p2ߘ�_sõ:���=�m��=������[݆�{�hG���Nf]r%v�~�sԡz��=�L�t�����y�?��_x��{0c�����ʫ/�Y�cΜ9��f� ��Ӯ��H�Ϝ�5t�J$P�N��O#�a�7���N9���>]�]Kנ�ˣ��?�|�>� ����V��K/�O�<r�{{Q%�_�`��o��g�3g� D�(�M�^1+����j��X�ч8�_����������c���Q�����ѵz-��r	���U�ն�-��E�����˯[o��N:�r
O͚��� �՜�"W� �b�B���#�h�v0�����]��p���Q-��PटJ 9�4Ƒ,��.;c�]w���nRo<���Jk2��فf浜�HTT�׵�8���Q�oH�L�Kus��LH�&�Fl�ʸ}��B��G"Q�RIDI$$c�2%� �o79��N��t2j�K�#��-+aʴ��"
!��j��-�Q�7"7�]�uߏ.:o�O<m�J0���ǆ��W�7^�i��x��6������r(��Ͼ�$�5ǐ���9�N��|W��_�֡�>�j*��6S��#ݧ�[�UQ��)�I���V$���q#b_���C.@���|��=BJV:�:��ݞ�+�I~����ƫ�D�>�l&���vU����5=��Z��շ�6P6��/Q6�Є��L�և��LV�w��쇽99V�YZ�"��$�0ٱ� �J"VE�Z��w��_|��)��u~�T}��p�嗉z���!�M?o�M7�
�.R����o�:3n��TC��W�Y��ڌH0�XH$+�y�1�M�:RIT(����k�QYۍ9�O�7E*�CG6	�?�Cgw�ߌ���Y�a舍�l���ӯ�q�������2�~(���?�!�fM>'��$��m[������(�28㲋9?�����N�����k�P��S��i���]tVt�#�h�{��½��_��ιs��Řz��2b#;V1"+����.��-6�GN>/��2���G0o�<�U7&���7��+�<��;��x�����<�7ވU�"u�/�WO1j�磝����<b2\���Kx�����;bD��kjR�!�ڷ�~��ē�8]�N??�,L�|��~{,^�uM���Zӆ;���[f�(צ�L�7+W�@"^���(��`U�j\4{Bu1���k<r�ø��_�e�P���\x��>}:�l�=�!�F[6}���ՙ�a��v����TħO�^{5�օ�8�JAnh��Ę�*H���Ҥm���&N����F�`�������~�����b�u�K��E��b��?��k_�Պ�lT�9t��ns9U�s)c ݗB8L�zH�,����=b�z�tc�Lg����R��%-H�x榑�gm�0��h��$���lo?ɧ%�H�.g�@(�N_�M6ƣ���㋿�0$���ק����I��u����̓�� ��-��o���t�1�
[&��A��IqF�Z+f��
�Y�cbfX}JD�Q�o�����%!ߏ �%�y��8�/G__
mmm�Ց��	�� �7rm
�*F���Y�ܺz{��?�����TbAAg�
t�l1��"�nhĎ����o�=�]3f��W^���G��V�Uc�޾r%��Q�c� J�F��\��������^�z�6Ǒ���>,_���#G�Ĕ�X��
���(����e�*�}έ���1}��XZJcYo���+�h��zc����d�j�}�y(�CX��ɫ��͊��,�;�|��>mԢ
���g�8�4��9~c���cQD���E�	.�u�}���蟟!�Wo>�h��;λ�O9Cw�}�8HM��E�G�<�V����PLe���/0t�(�=�r�畧��i�~�Ą1��1A�d���=�Z�}��6D��щ���g|��b$�Y9&M�):�PD7��ps�^����?�|"��^���˘;or������1�z��l�I8���������Ϝ��Dk:�1��	sgݢ�m��K���/�N��:
�4��"x��1�e0�>�0tp�uw�V�x����;n�]�U>�O�S/�cƏWR���|��r9�}�{'�`άE�J�F��H]=
�/�ɧO���߉!#�c��`�ܹ������}3���.�~���N��s�^��F6�g��C�u�<���?p�eS1��C�)�A�W}a�KU�D5��ɧh �=�oEK��`������>�$���UQ{8h��Ƃ:�`���X�\~�!�deo�5Y�U�U�V�����ܤ~nG[;*D���\�9i9���ժ�S�7���>�m[-��|!+oI��[� �\��W3TleZ����G����%��M8V�Щ�@�.�L�˿!��������e}�%�纡���;��k/l��\4�;���C2YD��`�lңyǑ��*���0*�簗�8�-I2�M�B�8Y��%��y����P�1�k4������i7��)��i?%t������P��y�f�I��� '�*�$a���պr�,�����2�0�J���F�����e��w�EYbU(�ݮ�[y8���Z�s���ϸ�QaMWb�:�Y���y'֬^�h4,��cF���_ś/������1�Ƣ�R@)`���8�`l��<�U��P���އB2�K/�X����梔�������kP������P���`-��u&m�5<�P,�hG%B�\����7��|ם{�̹��-�a?�P��C�Z�8�H?���C���H��p#�}�M\:}��z+%t���ы�SN��S/F�6�ʛw�)ga��1����2]���CH�=ě��^;�W{�������"��t���'����E�c�L�2{6��ӓ�P���~�W�r�J�鉧0q��0�ι���w��>|����x�ч��_�ǝwމbcT�tr���pu�E�q��p�٧b������ᶻ��R�Y9���K>����p鴫���AO�L/�1�5�oo��8~r��
�������*x�o���o�=��A͸h�%�}�=q�q�k�]��p�_}�����~,��\9�
<��?�fk�C+�_�iӧ��W���#�{�M�{�=�a�Mj�T�*�4���7����}�!R'p��t�OO����}q��/��t�/�I]�xÔe������a?Đ��qô��Ic+��┳�P-#�"��[�X[�FM���fߢk(�������DoG����k���x)�a5�!��6�6!� ݗ��R#H>�����k������f�7mX�f��ۧ
Ŝ1��kژ�*�ݿe�a/�̩�&�ӎڔo��^���Ő
y���x❷�����c�נ�Bf}>��͹����[F��nړwߋa�<��,��^�&�9�	���ֲ��l�d]p��L�[aP��X*9�W�\��Ҝ�SC�
fb(�L#4#��������5x'� j��ѣ�{�9�pmV��zFR��8vB���R��-�﮲����ޯ�!p�5{������\
b�?�M&��~|:�eA��^�+������V[��=�bA쌕��D)������7p��P��еj-�q.��d�a�>������0玡��Q/��@��c.2흸�+P�"=��0k�-����ixd�f
i�&�q͕Ӱ�{b�@O!�<=�@!�ŠP���Y��D����&ٍR��hT���n����,�F�F�Kp˵׉�:n�$�v����c���b�//�OO�	6�m�fR���[���.��|&�M:!��r�<���<�����⩨5RU�>]���_����DDc�6i��=��?(����iW�ʛnPu���gb��A8�����k/�7�t�!��.]�P�}�9�X����{��w?�o���e%M��~��㟘u�ld)Ų6��<�5���p�u31f����S@�h>XE>�EfM'�}���.�l*|QϿ������SO=;m�����+W�����n;}|��e�o��>��jD�>�p��.,^�5���FL�|V��]s�z�L��F����v��D�������������ƛ8��#q��NT���0��11�CC)'�-Y��b�p;���l̽�6x�z����I)�)�c+Q�R0��˶������sPJ���e飑;�v�$G�Q_�)_aI#��y%��ƌ�hƾ�)�!a��9��\�d'KIa5�DGز�k�Cwo��.7�������MS�p:jMcp����L��&dT�92��H����t��MF|����\����S_�!�~ǝ}��W����^0b�Z,z�qJ��"����M����e�s���CZq�-�dA�U��cA���ͭh�5"�*>��V'{�W��h�P����6ea72hS��8gn!ƣ����c� J�8.D7u�v}y���`A֪��-H;�����,�|���S/�]�|K6���K]`�(v��B�p���D�bK_��)�t�8\|��H�Ȅ������V������z{�)̻k.
� >^��x�#���[���D�WE��`P��`�C���B��(�c.z��p�UW�������_����ǡ�'VhoO
��!�N!����_b֬Y�~�D�C�s�(�`r@�?�BW~u�%�9�z����-T�&��D��J��;�y�5�c�]p������|G���pn�z9N9�Dl��V�m����0���p�%�T!�5k��������|�M��v�T���)�����TM-^�!n�z���:�;��Eem/�]�K�e�E�/��{���[oBcSf]~�6�S�����^Ɉ����G����6��oӌڟ�3՘��,�c�~���܎$=78�!��3z���*f;�AMX��%MN �,p�7�5�@�=?n�!�*/"�h��w6�GCOьk��3��W���P*#��b�ݾ�SN�l�= �y�m<��o1hP���D8���/��
8�Hl����z)�y�o8�4
�<
ZeF>ɞ��̳j]457`�=���UϏ!c7F �B��E���s1�WF}&���
%�a���Ct�p�r�t40xfs���.hvNb4C��f���r�0z���73g"י�Іf�{a���(��q,���C��^��{��9��$f�W���7+��<��j<�G�Y��5Gx�����	XnKt���PX[�u-M�f�n|o�ԓT�5���|cq�Ģ����4���,�O�����x��J����&z:����-Z{ӈ�3���p��a���.S�C�2D|U��P���~)�C����FU7$Cp���}�N'�,�e�9F3|�y�z��"g,;;�P2��r�&��WKhilBKK3���/_�o��M�\֌d/kn�_�:D1�iX������#��C�Ǹ3qY�v���ڀ��s.v:�L�7:S)|4>��V�y�dt��
@Ut���J����S�_/�W]=ސ&,��B<}���	��A|��&�&{Q2Аm�.|h���z�.Y��n��ե������_ߋ�?;���EG{;��,�}��x��g��ɧ`��7���0R��Y�ҥ��G��WL9S�:��
�r�igP���m�>L�z�2I,|�,x�-\=�J�uwb���kq�ϧ`��G�;�q#R�>�{���e�]���J�ܖ[n��#G��g�!)�ɓO��;n���_����9���R���%�q�����nƐMGc���x��?��e�FX���P�˝���B�Ǉ��!'�@�C5W���xB��=C��t䏰��{�����W��A,�49�L_~񹒵���]ɬLQX	">��ip$�ʅ�"V2m.@$A��V%x�FC/m��!i���"b��̈|��	�S.ߤ%!�v2�\"P��c�j�ːDӂ�%$'���2BYZ[P��+��|H��WP����X��:
�Ţh�f�5� �a�f��w�@6Ӈ�߇�D�l�^�#F#�77�=߇=?��G��_߅T{14xq�pt����P�W1n��FC�U�Wh�bܼH^��������U�ֿ�UW�u=�j�k9���6vc%6DW<���I���ZS�e%����xE�YQ�(Eb�5&0j�=��d�=^_���3�w���k�hW�;�Ww`�#�EKw�4��X?���e���������W_�}Z��b��W '\(�4�����̓@W]�72j������!��1�0��"x��*|=�L;l�K#t/W���+B���P�*ۛԢ�ОY�l.e�A� ��yU��f�k��q�C(�!��H�D����]���Q*����q?Ǝ'�]!?��XJE��ɧ��������_�<�O>\�7�|�-Ķ[n��N��|(�E�>V�5k�l����ݝ�#hnl�Ǫ��� �� ��2���cX��b\u�h��)�������C�=(}丱�� ���/��Ӊ�:��J�� Ƭ0%*��e�j��($S�/��Ӑ�S��^��-&��+/��+���g��WcȐ�J�������⫯���Ï�T�Ͼ���zW=���9��mfo�K�|%Rܸ����S[����.]�TbDh��!!�ٍj:��������֬Ų5kА�Ǥ1㔸udR�7R�R�)Io>�Ď_M�8�ɜn�$�c!�H�+R�PA��-9�Y)#4��4�z{2�,$W� ��f������"\
�1x1��SFO.D4��`�����Rĵb�]�m�q�(9[��"�i-��uN�dZ:�"�1Mdʜe�7�MCJģ�o�T9%���)��@���ҕ�	�ѧ����1$݇A>��i%,9��d�h�c�ؑH��2��e9,>�����k��~�cԖ�b��Y�K�1,ր�/,8�t�P�E9��獕��~��tM���
~v(����!�X�6��~f_��[�1�6�`�=�)?�^��O��<�Oӭ,�!� YE���v8��	���Z���o݃�mi������=Զ�ՍۺU�6v� N�-9A�jv��\���W�d-#�Ǌ�(HsJ�%E3S��*�C���@S]=���2L.���.x�qtgR�"�#�yQZ�ꂛ2��r�~M/�b
/�g�W�N��@#=��2q��eik���;tA�\4����@O�\cm�����T�Ëb˓N���L�ھ.U�QT�~����Ïau{�,?{M�m�9��kO��N��rٲ�����_L9��o�&+���$T��r�k �l	�� +�,ž��ޘ_��h�"��ʥ+��?�G��W�vͱ8�<�h�� �
���f=W�v��Cs$��_|I�(�Iҩ��I,nV!/,ÍA���i�<CH�u!!f�ՠ�/���D�*��%ʰѰFt��}(�ۼ�*�eoϏ��fU�4���K
v�����Yd9,��W��0x��Q�2>_B0��W@	$�Ǆ���дa��&��$y'X����zx�Ԅ�23�	��2�I���]� LN@0D[�ZD"�F] ?���{1h��b��:�C�\�TZ�EE�3-7�!��xŬl*�L�}�tH�4� 헽M>'���`~�
�ndL6�E�!�&���$7�< ����:�"ԡ�p,��7�y�����nE1�B�.�B�����77�����,O������ս�w�=����m\�r/H� �H@EMԨ1*��5F^0"֧����Ɔ�ذ�D)i­��3s��]_��s�}��Q�>��{u��s����{����[k}����/�������,Am���a�Lo�[��    IDATN�G����)��ASGeZ銤5��]�����Mѵ�{~�5l!�����e�to�ҁ�J�����[��)V�¼�}�7Hq�Wy����
4?6��X����۵�]'_q���P1�����o9��ދ����x��_Ax����DN"=�F�d=3xO����PI�3gP<��)��X�����X��vBLP�����7L*�PYI�1�8�eN*�r&J���|p�WC�W]*-� ��l���w���KZX���>�$���V��eO�[��^��F�Xӕ��T,�e y@���4�c����/��^�Z�}��b!���M;�1����/���Y�J%�a<�D~` mZ��2��o��?W����.U�Ŏ�$EA�6�#���.L����#�MV�Q���&�~7YvMf34���9��d�%E�XŚ¥j�L�)!�=e��]"����%d�gקrϗz�#�Sِ�7*{,Z� ��ʦ]D*�Ѭ6�gG;��h��_ �}^ZdQ����U@˕:�� �L��1�Ř@(�3�d$���B Ъ� �1����Q'�"V��p�QY�E�����
�UG��`5(�Ȫ�TYE��B$���"� ͓�,�.{���ȥS<��+/��B���@VUU�kMe�h��G�`�4(��Fh��]Hތ-eƭ�G&�Rf��O��]�N��=g
&$M�E	R��R�q�R%�H�!��.�P���sP�i��e�"ЖE�d`����{n����X]�����:������F��2E��������r8]���'�H6&����F��xI�A4���=�j�m�U�����I���hU~��h���L�$�prɒ8T�#""���M`3����S��<�N����>���S��~�2qy�+'7<|��Z�@���%�{[���^fS�ʞc^*��$�@�c7o��w���.3=���(�1m��1f8C�h�$�X�����長=YH��3��ȧ�#hP&�uki�?���A��ْ<�L	z��l[�70Ϭ���-�}���#��&�@u��,:���`]��췼;_�j�4���ѬV�Wu��3mJ,��z�=c��k:&��iH2�o[����%mۻ鰴���iw s{ ��g��	Śt�U�o�=oFP(����ⳬ�+�o� @ ���is��z��P,ZM '�k�g�F7�P &�������$�b��`���*�؍6��B���z���IĞˬޜ$�]��iS���X����J��J��
UEz�>"Ɛ`�q��wĚ�Tf�r�T��^y�z����� �٬�n(����N�C�|������|~q���l�0<�c1���ȡYh���ο�
&����d�ɝۙ�u�o���Y眅v��G~��t�Hex\�i�:g�4�E%W�1��cP�Ay��h���X���=�L��듫��25�j��Ԟ�5I����
���4�f�-g���dP`6��4�Іb�Zc�6+�J�%�!T;-(�0�F��������"�����b� �X�x�<�yA3�=_���w��Y.q���-y��D0�<��-8�ռ���Ͻ�6�3|o���o���^��0W��Ƽ*�D`EGxd�� ׫8ܨ�r�?���#���rF�~�O�%�,|d�<��o0��&R&B�dP���E����t�lE�����d[������@E J!i97[������A��C7�B��`�R�D��V����L���D Fc8����..�_ϙ�(k�&�,�oԴo$1��:�Aq�6
���E�[Z�q��JXUu���|�k �j��B��%QYТz�`� ]X��J�=�*��P�F`G�u�-�~/�3H��b�x�-
L�&!���5����fD�L��Z��n54�lU�<"E�>d\!�hY��4ZMvcJE��K*��`J���CA���Z�Ȥ%"%�~4�%OUL"�f�2X����v��e��ӹ�J&� �A�]S�m�#�3��=1TEO�V*qy��L�wXW�"K:f�znF�X���[�C)��/����N$a0�M�=�dtZM�ʛ<~���)眃�o�����'aey=�&�Fp��`}}���6�r�8��s�%����p��)��s*��ɐbb|���6��� aWF<�8ӂ��K+�sh�@�L�5����!�U��*(���~�H�D���:ӳodm�R/��#��*�-�q��q�>�z�yY*��u=O[��¯
h�Kl*��2I��,U��6��MA[r!u�<m7���o ��3e�T�m�[Ǣp�6��Dϓ�+_��T����i��`K�x��xY)�gz�7-)���g^�k\��K�Û~ت����b�!�-�֢|���1Z((:��������p��2����~�e}��_#���rV��G7|FXZ|�>W�c��-�7s�B��hB_Dק�%Y|�Oe�^ɖOR�ޥ�eOZ��T�镉_������9�QH�L�Q"��;&�(��U��wtn�J�]O��{��@ �62&'���ID�27*���XdR�Jt�j�ˠ\�k{��ҵB���w�0<#lrF���	*A�zv^t��c/��L�mv�`]�IF��.g�6��:Ěf�o�v��rY��n�M��iq�jԡ��Q'Z$�Bp�i�����ǰ���i���d�2��AJ�]*%�� ���/R #p��1iRs�ot��"�E.� �8�4�=�|$]�Q�����\dI���(�A��!M�TZ'�6�;�H��V��>o2�����*/�h�� � � ;�L���K�޸I����M�K�--#��2Kx��	IS�N=�L���Z.����`͢+Đ�>+U,R;�
r'�������Y(`����|X��g�}��چť%��/"�� ?��^�#��
�d
�O�����F�BA�w�\T��]?�J��Ü�.9�k�|f�Y�{(��U�#A������Hz�T}�Y�SaK�6)CQ?��"�g����(h�._�9t��ػ�GDl�3V j>)�F_�9���~t:�5�g��M� V5K��ˤEAcҖ���F\S�9���")HZ�
d�ж�y��L�����į��/ɺ��T����5�$G�'B��}�z��ጹ�4D��M�=
½���=?cΔ{���t-�hܐb��	-}Ӣ.a�w0�B�6Q���_./~����e��G�_�@x�	q�7��uum��O	Dp���p����A�O"��A�ʠ�!cn���;[=�Jlc2�>� �⼬����0ɽ�$��ްt�C�ӣ��g�tä��Qu*��l¼q�D�#~=�}M�b��҃Lh?ۭ���g{e�C��e�wY��7���(���A���q�D2��jo��W�$ ����E�,�/�6�N��ϧJ@��ɫpZk�dN�s��-*��u]"^Q;���HjF:��
M�<SEM����J<�CuZ$�fD�,��]���r���8H2��H�c~i���t���9�4��e�ih~��Qo6091� ����:��r�,;3�������4��Hq���>�2h�����L���
W3�� ����7��T��������|~��Alh2� r�ǚ%�O��G�U1�����Ϣ��|����rj ��I,�/acm�l
�c�[X���,+N=�ܧ1����A:���?�67��cرc'��:f�����[Nm�H"	5���s$E�,�)Gj���6](UxdV�"���xcU��ǁF^z�"|e�Fi�ז�S����`eb�y��r���L�5��X�<DF�s��稂E-"�ϗ��� K�6�/Y	+��� �"(���=����P�Z�{-$�~��K��j�L�� ��Ó�=ZM��W��j��J�t���"g����(�jk��q#/��t	�gҪ�s�T�\skk8���pjx����>����}���[Ύ[�������;�c������Ј]l�������8��y�����	��Ѝ�I
T��<�s��AL��=�s���w��2]�^+m��7ç�i�.H"��E�5�n|���;[�#v&}Q鳷�����n��<�g5Hc5[-��bL�����#���&&p��}:L��L��"�E%�ރ+ .��� �ǫz L}l����bF-�X(K�׻#�T�q�i0q͆$:(��	ZGAP";n�&"����N��6�R/��iC&@��2��4�0m�>�g�Pi�Y��A��4�q$�K%�HEh�Z�U�|L�#�lM7�0� �E����l4���΀H�[�ݒ�'-�li�~�c��)ӥ� v3g,C�R��赔�6��E^�PfJ�Y�F�c �k(f�+]c��Q"ؑ�^ 27������������`�P@�TE"��`������P$�SO��~�߿�&����u Uh~z����0Z�O�>�`(�=|ݯ�X�g����p$�-M��Sl��e���
��86k-�K�$�� �H�}��7�c��q!-H�Ұd���l���.��|]̱uݵ:���ܐ(:MIrR��ȥ���ŕ��#�;-�~)�=�2%�� �,A��~?�7u�Lt�k[Ԅ��y�Ju� �wK���m;c�a�X���:���m��yD���$I�>AX����(�dY�-���8a6�j�$��DEf4l�C�M�q%tI꺢課L���́h*�i���N��lNX����;]���׍��+5C�]�/�'��[?�l툂�Ǝ��[;F�o�tC��K��K_��?Hs�'����o��O�}�?|ߞd�G����B�6��(ϱ��G�ᓲWr޺aӊ�@�s1�{�����j�r����T�Nz��-�7e,�N+j�L������~Μ{%7���Ho�Q	8.1z%p����i�6[[���x�B$b�`t�
���cA�*�ذMz�o/<�������:�\�ܝF���J��E�&��n��DA�|� �Jl\Q��ҍ��"��ҙH�m�5�-On���M�����$�&b� ��Q�X�p��d��V�J�2�f�L4�KS���@��2_�L<��q���%t-����3�,yAB:��t��!*M'#1��7Q#W&Mc�"E���9Vda�|	�	4�u$�I�K�q4@����4�'�s5eey�ߛL�8�_\�:��������(;��K�̢����}�61ɋ����� 2�X��q��4�9.AWu��ڱ�v�b���}���������{=ƇG0��"
��1�)~�p���p*=��?��P�]���L.7�Q1�+7˲KTQwt�~�Tm:�N?l	B+62p�?�_�˛�;�p�Z0���%�-H��AI�\c� 	����ܕe��(rC��YQ ��|�����_��>���sa������������v�mc"Ro"H����|E�'�ȶ̊zJ2�.�r�<V1׆{`遲yT�n�L!�#bS٘����4@=Hۅ�$
O}��xt\�q3~G	�q��#Ks�T*��K.*Cbt.mњ�G�i�R	����/��=�?\i6WQlɚڤ,#��-V�e��5]_ ��ӵEö�2eAQlEtlA*ɪ֚<y�����j�S�����Ӹ�*�H<�TK%)�jIm�_%+�����*�.�K�ӓ�e���AM��b��������tU�_U�IHą
��r�ReiK�?ȳ����Fc2���M�e�<���*�T��/��U&�P�H@H�ٕ�%�a�fT�*�b��x,��[Z���� ��2����2`���D"�TU�G��{�����T"��0����kgϭf�Y�t���y���^RfI�\�2����@ a_����<����116�c��5>ީ�	�Ӄ �2�������|��K��~�]?c����1�-9�����`.�=�X"
)���?�)��ɚ� ��,X�ւM�@RF����������;�z����-}����{�7{ˍ�����~���aw8mm����*�j���l�@�f�V��>��E�J�Le$�${=*�2'���� I���9u�~�aSK	x=fz���z7��-��ָ@o��7�C��-�]��`8��2:� ��麖e;�$��(Ɇ�ڮ�(�5٧��l���b:�{��??�;���w�o�[~�O1�~�@��va:�#Yd1�WZ�&����4���G����بV�ĮC$T��b�MZ��x��@w�N�7���ԭ#c ����`}f��Hm*�L`uy��2�N0`��y��������y�;?8 ��s/���I�������5^��xQ@�,T6��,� �T�N�R\B�s���x�睩�Lf�4G�ľ]XZ��0������ �ϭ,axp	=�~n4��\pj�:~q��|�?�)Oa�}�ދ�����8�N������옘B��D"Cj0��w':���u8��H �ۤ��{�&1�.	����<��K���'�w�N����8����ܛ�)�zh��ˏ<��	=4�7��SX�Ւ�n'hY�.8�$dF�2�u][�����!
%EUT�m7ֵ�ךLZ�WdK�܎�C�����"5J���RŔ�|H;K�$��rMt�2 �b��:������i� R]݆�	�u[�C4�/I�,;�NgI���󮺊�O���^�Ɠ�s�]YM	E�\L��ಒ�I�مc����E<GX0�������[3��2_R���U0X1L�d�'�I�,�ăA�W�5*El���OҠ�g�������R�E�F)+�T*����-S������;�G�F�`*9G�t�-�/0Si�@���i��J��;��п�=��i���ظ�����/=�YL����<����&�FX�уx���Ӈ���3`H"x�a���ٻ�+5w�y'b��6��p`��h5�H���d(�B&5�<7����6��w�I���$q$H�)�1���E_��kO����������?=R�``<7X�%��v��mG�(,��*���8��8�&�ڊ���h%���Uoq��J�M�t*��aY�ՕL]w������T�珂�c'���]F� &��N�ŜȒ�o�����W�[�r�[�::{��̵�XJ�XQ�֬�C�r�H=0���U��&ቨ?� J�!�|+�JfJS�+���kP�����ts��n���R�84����g��D
cc죺�.��S	�L,e�Tq���gN?"GQϝ�T��2�Nd&b�{���n�_C���1�[a�$=�m�S
 ���Yb��`,�%p٨6�K*�-!��p�:��m�A�����y���8����q�6Z��ln �����t6���裏2���e"!�H��P�P�ѡ�b���_U9��i~�ܰx����Q���x��w�s�����#p�F�����߭��|�U��}���)b���3�:�������Rf����Ag�"�F~�<���[i�f�}�Σ5R�"ml�T�4�.��yҐ4���H�#(���^m@�H&��Dkk<�J�m&����g���R�J%b��
� �~R��C`HYj�VA8�e��	�s� ���etʄ	�)3�Yg"X�V�ZF�Q���0K3��H�b�%xp��Y������0�����E��B��=�b@ߨ�����hu�	��&�qp�+_�#��C�g�dIYm�����"� ��p�mO,����P	���;��J8Z{�On�����-�#��.}����'�_������#����i@�m4�.,udf��憉J��0 �9͇Z]�_��/Hn�"KZ�.�n��AC,l��,h<.��4��.���_C*G����J�D"���)X�XB�V�@<�D8�@K%dQ������w�^+��@��NY9\�Vf���PVHs���t���옶��x�+��	�	�����pI�+�sH�#Ȥ��Y[es	Ø�����q����"�N"�J��G�������6����n�173�SW<[�    IDATO��s�K�T	uҪGx��z��x�Y�ԇ� �i�]�%�f�3cR��H��x4��c���E7�z���S������������%_޳��Y�p�4��ζHQu�	=��a�!����@�xW*%(d���G�4�E�Y$٧��3	���'�c�݆�m@�N5�M�6L.��EQ��Tʛ����$X������T`z-)��)��l��[tL�J&x	L�wʖ)+��.�o���^ʦI���P���3�o��afa�G��g�S���Ӈ�ǡG"X\^�)�ͯ� ���e��x>��Çcjl>I���<��).�g��dp�Q4�n҉&�e �SmduA8�
�&��مԛ�F8�Հ�|�������G?�������{N�|��Kޔ[ݼVm4�v:��dJC�`~�O��J(nnbll�A��͎*azi	~��ZG�D�]b�;h���Bb&;u�`��z�]��d���1	�	�Q.�xN�p��|H$"(�l��Q�]_I*	hQK��|��bs9���k�ʹ�T���2[z���0�+�.�-g�++�=�3OOOcdh�"cyqɛ`�Z������H�����<�Gỷ��3�4�f����0t�6l�-�e`(�D�kȇ�L�"���v��۠�ᡥ��j���#v��`�@IDcq��%T���F��mN�"Y�`�X{я�̝P'`g����J��G���7�>��Fڶ����lM5�{ր��D|�H.��:��$Oh��X��$�~�eMa��]4,��#�4�nut$lR�YS�R�VHu���D8�@�RF�VD8("�#
aua�gj��L@I༥`E�Oԫ���_���)�����>�zI�*�2�SI�2R"XQOwey����:tÃ��󼺸̀����Y�CO��`�p�ӟ
1�y��z	ۧv�[nf7�X(�}O9ӵ��u:|�����ý?�z���P��{��!��rX�D�woǣ��m/��Wbdl�����YD��	juH�T���դiOFG�QG����큾H���e�{}�}����z���>��{��l�Ŷv�뻩I8��g��Q����{�g��|*�luÉ��kP*��H�.,���t�مK�A�b�U`v �-��*���h(��"��Bl<r���M���d$�Y.�����Ҩe��;�m4��hO ��`LޭT�ެ��$Mlfc"[�-�x�V�8fffx�x3��Gc���X^X�)���q��?'��r,���A�/�%��Nq�|�#������J��C�{�17��x:��Ї��?ƾ�Q8��
�h�TbA84>��ً��w2cp*U��u�C��>�Jb���(C'�˂l;�EMEE5�.y�A��=����0}�=���.?��z�w�����Ǥ �]"�ܷՄJ��ޅ�?�B8�+��`,���ZD���uH�&t�0m#I\��W���{7�C��]w�y~|�yl��W\����pE�<�b�Q����&�sP����ܣ�,uK�y�,E�E���,e�D�"��̘��N޼������\�`4��do.wc�+E����#G�F����~.5����6 �#��?C�{5�,P�_��_�6�J �y�+�����W!�}�RQ|��������������r��8-;�T(��6���I�O��ɗ>�� n��]�Q�_�u'R����<r���uh"��mC4D�xº�o�}c�'~��q�D����W�ߑc�������h6��袆����Q�?�d<T\�K_�z��zP���-ec��b	�m4!֛,����������_�*\����Vo��mxǛ/ǳ�;>�9x�_��������u;~���cG@����Vc��̕��4�K�J�J Jĥ-��f��L���4�C:��0g�s�\�%w"�l��E�M�N����x{�h�Ã��>���?���u�ZZ.yj������;qΙO��>�wx�{ޅ��8�9��w��e<���ͯ=����ｨ?� ���bO6��'�R��v�_|�L�=r�o|��a��ގ�mb��7,�]>W@�$7�M��	��Cj��u��
�zV�X�/�m�#p,#��c������肋�M��y� X�SF2ZR �D���s�C"����c �DP�����O[[Ǹ�G�e@�� _U�B�Ɗ,�ɯNzџ���o�]w߅W�
��G?�s�~2�J����}��@h��ޏ�c�bX�QYY���H<�lf��R�M=�d"��UT��7L�"`]^^f�%y�����|���㱢��Q� �&�ʜ�\�N$9N��s(�յe�2�D☟[�$����B3����ԩ{��w��{�����=8�%/� \���s5����ܑCx��ތ�[���?cG:��_���4ʰ�M�p�E��2��c��!�0�"6Z�F��'��R�FL��촡h2\�AD�L�����w_.���s�\]�y����X��'d~��w<k���s���٫�E%W��k'v�����]w��QAm� ��")m��D8�������laD lXX.\Eæ�`�V�Y�r*^����������=oA8G0��G��>��66����W�-^��y�uؗ� "�˨��^ER��j�j���x�4���6/�J��#<7�H"��~�/,/yR��Ø���L��'���9O0 �"Q�󮒜�"q�yqn� #<2
�8�͗����5���>����>u-r'����K^�r��B�h6p�>���A4� �������m��N����N�U[��W��h8��g� %�pva��f��Btlv���!yϦ,��ٗ��q��?���'b��`E����?�<�WW�9����N���6L�F����A�;&���i?�4|�3_��n��3���.UYr����}��MDA��T�t�;�T�r��ȏ����׾�-�"����s~�~�Z��ꏣ���X_���g=��}?��W��ژ�d�'�ʍU�n�#�!���h5�iԡ(����Q���E����7
bia���*W�+���4L�/�������.u,���*!?±�f�  ��0#�>���9��*����`$����1FNE��� d�����v�t�0����&FG�p�zF��8���7��?�9lW�Զ	.s9xk�"Ƨ&q�]���_AJ=V���q�d�hYh�2������_��?���������������"��w����n�E��@��0	-IF���K/��{߄��|�?��FT�9ˊ��ػ{�G�p�u_�h 
��AD$�v	�|�{�ۀd�w1��p��߇��?�,o���n���>g�q��u��э����^G"�b7#bR��V:�@>�B�X@�Z�2r�Z�K������d*��K��[�����3�0�x)k&�**;�E_*��ꢷ�@��#�N����EV��!,�,#	#�L�Z���o4�0��H0�j���K���:{U@>����i�� ����� �H�^�`bb�R����J�趚���뫈�|�%m�]$�-Y�z��>�7%��~Y���#p�F��'�7���'����}�?�ᾜ�f�5E]AFݰ1y�S1����� ��2ґ8�V�e�\+��眃�d���Oa<�E�X�D>���E�ۧA�B0H5�AC(X/���napp�R�Nu��X<�`""	H�:�j6�E�d�Ґ�g�F����UL�N�X.�o�?�V�}H'�<�����*����<�x	���r�?O>��d���g��`qqR�J�qdv	�?�L6����Sq��8sΤ�X^]�����ή���#���b�&&��0���r�-U�%H�~V��F��@<������4	N��X�G#ҞǴ-�	��0t�����7fB/x��:�/�G�8�@x��/��+�.�]u�޹�w�U�b�a�2\Q�e(�&�� ����5�%�|m�C~.����z��h8�,`2`�YB�Ղ(�`�Md�I~����-���]oA�ƒ�Mۀ+;P�(����|��-��y]���@�TF�����ɣY+�y)�%�2�Q����	 	�i�7����iD����VD�A�!�49��Y֋p�t�+s�QO�0?�
�/�\&�E��l�޵��i�dsC�?sRTg���T`umD2l�
�
�0��V ��([&d݇N��T4�T$����m
X�(��0�s
Ӈe,�]��.��!��i(&��w�kR/y�g���#pF��'�����'���x�ޕ�~p��c�o�8@ǲ!�
�fN,��w(D�|>X���������{�R�G�T������\8&d���L��Vˁ K�ަՆ�`����iu��u��r���6�8餓�,�nP�8ŀI�A46txڛ�%�F�~%EfP%�&��t� y<� o�{	l��l��\�2q�/����G1��ѕ1><�#�#��AUE�K���~u�1�3a��47ꈆ�b8p� B� "���:��p�(q&�������	f�������(�,�m�}{�]Շ�����Xp�+^�K��UkO�,迣��#}�=>���^���-�x�ꭷ�4)��ڦ��с-:�B�i4ȱ�I��&��V�\�Y�$T���0l��� N�\H� �aA�}0m�&²�* ��>]C��r�(���D�� ��a�MOr�l�gy�� �����2o�܆"���m��YL�aa�T����o��������
###��(��C^�����Yf�\&���9.;����r	��b|h���j#;����Z��G1sd�H�t3�KȦr��ϭ,����bmy��D(��
�0<��(�h�6�ut�4��F>ׅ"
0M��m;�Ϗn.�}��l���-�S���~�Y��{�B�����G��j��nx4լBm���
�l�,�ir�*)
�6Ee�:���4�uĂa�Ri��Z�k���`�m8ee!�&`:6�ܶ��e@Su؎�N���?�V�	[�أ�ӵ!�B�������d�^���ju��c���(o�P�,z��yD�QDBQRʄilh�\�,��w�dMs����	o/KQr�h6��Ʊ���f���W6�"�� +ҹV��0�F�9�/�� ����3y�&��կF`()L2�%2O�IV�I�0�}-��z��.����Fr��#]a[I�ʂ( ����Lᔗ�|8q�e��W�я�	�>�_Z��x6���w�_W��*�v����f�_	��Ȱd�(��Xl�G,_��);k4����	MV`;&�{]����2 C���D��@���v��	`M�m@��БE�>� �m`$����
�&wlGq��f�#�U˨�Kqju���;�������2^Z ��2eؔ�r�l"�����<0����J����A���A�ǁ�ڢ���gU( ���&��Dz�e(-MA8����y��L�(,�@����,i@��!H:,I�����Ž��\��F�	?}�쇻���@ "UD	��UdH�M������q�}���'~��я���>��C/�q�/|A����n��eD�1��hD]�S5= Gձ�h����Lv��>��	����d�Zg�)MA$#Mǆ��X�#ȥQ�Ԇ�ɐ 0n�P$�"sF�����h�L�F�r�w�EauM��h2�f��r����I�k�Je��XXY���Ȧ��L*5S�K�-/�x��7�T.3���E�<04�j��Bi���X���j
l^p��:�|'?����i�	,�,b��a&�`bw.=���K�x�QtV����b�\@��B��J�It$eǄ�	����)���⶯}GD�0Y�$$p,����Bp�#�@��O�w�5����2���#p�"��c��������g�W�vL�#�����3����� �u!X$Yh:�9@L�Yԁ�������[�CVP��ܖ�E׬�� ڕ|���/�k��e�	Q�a�hh$E�\�"�(ؖ�ba�UF:�C�Z��f	;ƶ��@��� i =�2�ms����ES�K�*/e�[�;�`�5:���\��ިad ���3
:|CC8�qɕ�s�,/��o�)�H�ލk��VLN���^s�L��0�@E�{�Ʒ?�OSDL�2�YY�f����8�PKfkFO{�E;i�t:� ��o@sv�f88.$�#��ħ�8�df8�̹�8��~������O?�k����F���>7_p�C���S���w����UT]u������8�I
��g:.���$e��*��
��â��cc�S���/�c ��������]/~.`���Y\���Cca���U�|n��ǘ��t/��w��8���ӿ 	��<7��bpt�z���;ƧЪֱY, ?���*)T���r�n��֨syyk���w�|�lG��x;�&''Qk4xi��	T�K��lBF�ԝ8��d�����/a$��K��|�3��
��o{+���~� >�����7��L�[q���D,�=�Z�U��5���i{��x�����4�8������������ms^ _^�Y�M"�䧞u҇>t�	B��6}�������ܽ������HH
Z�.�`�BյQlT�]����?�/�{����_�a��Z)QF�kA6,﯉.|'M�+���F��¹{΂���5�������y8r�=��羈����~�#x�;��u���x��O�o3P.�S/�3i�Eem�5�����颰��]��Ѭ�Q�XGv(��b&[�'�U*h�Z\R�r2�,��4�0e��r���ccc��6j5l�چV������(oj"�Z~ ���h�@W�v��G�;^���a�TB[�pֳ�������~	�~�`ߋ��O���1鸘Jİ��K��u��������_��(b����(H
FCI�h�8�U��v�{#Z2\h�JKAۻ�٧���������S�����m�����7�����^�m9��W	�٬!0���9g�(��'F������߁�'������Mȭ��.NNd�)n"`�좕M⼿�G���? K����W�n��O�cصs
/}ۛ�W��x���Y��s���/5�nO��|<�Ig⃗]�ݩ8v����P,�al�8��76�8e�n4k��� 7���f�k!ˢY��R��Pe��Կ%V31��	x)�eQ�j���;�S��Z���P�J��r��q�Z�>��0]�'>�!���obci���Հ��[��?��j���wq�3/��矃O��2�R$��#X__E��A� ��|�ؿ��#@��M1_ Cz������?GX�aT�i$�����D�:��>��_zS�t�G�D�@xO�o���O(���\��.��R�4��lEF�4������g�'<�������;PX\CPձ{�4������7�m���6Жdl�ڑ8v>�B��̋`h�P]\ć��{v��k��+|�����{�� ����O~
�w����⚗��$b��QXA�YBf Ϟ���&��<�zK��񮖊pz�۪�Q�T��L�-b0����4NT�T�lE�e*9�L��m��+H���t��m���h��x�߈ǪTMg?����b��G�k>L��7�g��/��(x��;�_�����v�4�%�(��X.�P� 1���핸��[1=?����~�A$�L�Xy�!D\F��t0 ���H�YQ!�+<��R8��Ϲ��/zB'@���G��q�e�w��E���o�����l��D@.�R��A�v���ݻp�ŗ�?�9��J�&	h��n� u�;.GR SR��b�Nl�#�M��,���A�����׸�O_���z�u�x��㱄���    IDAT�݈�t��Q\}��kr/�����U��rl��P^Y���8�e���ݷ{�&f�g�%9������,���,,��ɼ`px����w||�j�����8+&&� "��+�������6�#�8Rk��?��1��������_��=g?	C���'>�O
*.��r��,/��$����$"a����e�P4��,#<�G~jS�����5�{�]�U�p660�h�ڲ�yjˆ��i7�5��W������cw���܏���@x�m|�[?N"P�����?z�҈��|�.l���Iп���*z6��� z� B>?:�6{����mv��F�Ttj(���߶���E[0ZH=�8���*� :<��}�K8��`}fl{csfmel۶�tl۶muұm۶m�c;wlc�y����O8��^��1��-�������3���l�j������7F����:�a�������V�ֺ,�`��3^[�T��]y�9Z�~1���ZS��Hɠ@-��=-Qf�o�x�gzY;gO��1q�oR;��##[��~�R�i�jDbI�*j��,��C-{��O�~�ҩJ��Ǚ;v���މ����Ppȁ:s��Ӝ�pT8����7v�ؑ2X*f�篟,�+!i�f�z��FV�<�(������];9[?y���x������]G��@����W�1��<{l��,��<�߽|��=���z0b�Hk�~z�G6���k�8	E�f=��_Шe7��4^�Jt5����1=�i�q���Xء\�����8A"A��j�j�1���vF4�>.I���l<�#ޓ>��1!�sF�� -��`��m�4	U����`��J.��f�t޲�e�vj�G/�F���Z�I8�%Z6�
��b쫦�v#���a�Tiȏ� .�j�&̘�:/߾BMl/�&=����m��X�ӎ	���5�wQ�B�+9�7Q"+̈́�pd{I��c�:�c�C�a�D��Q�n w}f#<	�_:��k�>NE��<�zn�	Z��n\��YX:��1O��i�>��z
��2(��T�b$�օ1��3i���|�Ci
���4!�������K�hVq��sl��K�(xZ�@&HxH��q��(`0a��1��g�ţU�U�M�*Q{<���T�G�p�1�<�Ħ3k}\�w�����dէ���+��emjJ/dq+������Ud�Z�7u��T���Õ���3����E��O�v������5'I4i�L���B1�6H�d�srr�%f7k*�aWR� [�o��s�H�z.rlܾ����\�����v��t:xF�a��T�|j@>e!�?�~Ϗ֛Z��gH"�.�i[*AT'���^�))�
LM&;��8J�K+"���5"tmn3�������ؓT�y�A�7�FH1�v���3q�3�lP_rG��Z�Ag0�&N��P���4g�GC���]�1�L*4��d���Op͒��d�ܚ*i F9%�+id����ƲS��`6�J����Rza���%>f��CU]K���;Ԧ@��4o�h��6|�l����cE���n����34p�����,x��lǒ�;�P�r`UZtU7�h�;�*Ep6
��2��+M
Q��x0sۮZ !�9k�}I�FQ��� �^�������p<ͧ��'Xq �˦��.��������aQ�)�`A��k��D�U�	�-6������_���ʲ ���c�_��qh�h��q��E�{�-�^��T�����:�dĢ-Q~��u��-s����I	�Xب�������`΃��nV$*�֩)*1�hΪ��FUٜg�����'E��8YIK���ߓ3'���I����u���3��G�x|��+��jn���	�����GBNs�؋\?�"1r렓;b�\L1Co=n-&{����%�w#��)��,uqԃ���?��ձ�/@��9��-��P��������ȄP���me(K,�nQ+ը�Cv]�h/���x��������՚n^�Qwҟ�=v��l��βp�d#�wl�0?_���X#�g���gb�GpS]��oك��fɧ�Ź#6�hqx�����]��*<]�ﰦ�\�
)G1I��{ǖ��z�M�����n����@�/������e�F�Eϩ�ˬ�/�q9�XU��Vs��<62S�.�i�.U�>]f��L�mq����YF��5Yb�ig��O�o��� �`���M@k"�㞈�7����X�7.�s���.���'��!b�o���舙#09o���9-�(& ��Y�U�G�b�m�vM���PY#$Y�z�`��!��x��J	/�N"��zw�M�!��t��XP��%�jgo���j�tS$�+�W�t�mW��N�ڴ�%����p1n��7yދ�@H�_�����%�2$�`��2���M����DZ�2�UR����Cc1�yW0S���­P^ib����@��Gnq���a��Aܕ<�_q��`.�N�@�T=<(c4T5�R:fhk'�twv�w�4ٱed�a��3�q�B�������ki�c0B<�э���k4H �݃O���5�o�y;�5����l�?xNSѻS�]7�dS�ZLt4�����gꑼك���?�9��g�䱱�bY��ؠ�hj]��ia?g��6ܶZ�\�K��Di�M�C��{/�$������d/~�u9a� ���Ү�����o�u"+�X�os�7/�m+�[�Ѩ��Zm��o��������b�s�Q�:�]3�%A�Dq��1�M�q/�r��U�P*{�H��u̧��KzrΆ"�	Ĕ"2�7����7�{j����[c��h�����m��"��b�3BB�C%ھ��i��lu�Z�x��[A<�&�Y�%���O{��m7�AON1 �Ph)Ǌ�7oy��o�o_��v���X�h�D��z��}�4JD��Icj�st5����}!6i�8Cن>E�m(f�M-����T'�N�(���������|�ȳ�,Ϟ����8~�U��Ld$dK`|>b�'�����mX��1����*��H����O���!�_���|}�f��/��+'�?Mf�">��`��W�P ���S�'���QH�%���,6f߻X$&�VF#Cwݎ��e��O�4Er\���?UW�wBR��*i��|�X;93�����(�`�R"\4�VPo�.�� cG�P�E� /9�Q���OÓI�9��+hv�8PV���^��p=���Z���(/1�t��it�׻R,�f�������(�>D���K�Oʇ�.]���$d: b�;&7���@9d&|���'>�nh��T���#ό-�L�z�&#�%mI�y Á�V�A�HK��%��i��1��aڿ���7�ڟ����1�}8��Ք�U��n7��@N�1�S�`�.ɪM��r�S�T��?�p.!G���`��e6�����VTA���Y��U/�@��_���oW�#-Rm�!����-��zo�y��	��Nڗ��ޫ���ʔr
��R�hml Ka�x�	2￉�
�g���S�E	�����rI��	w��9����6r�Mh��"A�c�s��}��`B]�]"����v��w�ꔟ0�������w��߃?��}��ݔ�m��wFf�?K������̙�T�L�oJMuCb�n��6+M�Q޶NH�m�6�� ��5��Q����.uB,�K��DO�i������BC`sA���O�tdg�<�F��d.����g�i^��h��e^D�VZ,�z�:2u�w�y K_�ƈ�(�,�'��R����E�:5������ڸ���q��An��
�85Oo�u�|��++�U��0 +��=�f�Q��_?�i�W���E����M�B>z�r���'�6�l_����O�y)6v��v���SU$�pw��LNN�?��xX���;�f!}��	r�����-T�u��t'/�9�\�K�}
����$EOW�A�C��|R,�܉��+_��� ������'!5��Gm����9�
\i�_�,s�yׁ9s��ӤkBs/������M1��X��V�85�D��
�m�Z��N���,�@����7�y_�?� �~�J`��T�X52obDp"ǑEqڳ蜛���0Y�"�d�R̛�����9調o�#U+�MZ�����>L�b U��7@�"[��������n��F�솤�ւ���jwh^�����U��_Ԉ�f�ǆ��&�����@�K{���?���x�*�Q��?�g��$�2��T�Fc����3{@F~��@�4ߕrL`�Ō/T���s�2 ��m�vr�@�w+�,��Q��������x��N	���/�����d �5f�>0IW_@<������+�8�)�����Q"ƍ�����%o���3	�<�M�fOO����;E�ǉ��!�'E���m�S������Y��\JV�Aze��*�lwF�ڮ��eޗ����OP��t��	4�/�e*G6`���j�9����RJi<!���?�ԉ4��d�����i�)��i��[")�[xv���;;��A���{JNz[��	e�-�}�c��(�<�;ڳ���g��wٹ��}Z�c��S_/Mgo�Nsq� �&9�A�؁� ���D�k*#+��/�vj{�:M����t�7B�㯼���p�J���錠D���%U		�qg��?HH닮��#��~���!�&��Xy�'���K�ts�
��\1x��z8B�<w�ۇu�&��P�)G����k�tß�#��~���5�E�UX��s��P�}niawB�i��W-�<����=7���Zݹ��B��"Aba�ZO��
���K z�J��묒�%�c6>�N4���J����U�	���3�3:����5&�����y/w� ��SOW1�����4�<eyjT���(�����cܛ��\���<��Zf�X� ܾO�ڟ�:&ל�^��پ��4�Irq�\Q� ����V��%���9�ISI�f\�{��w����Z���r"���\�o0���O�Q���q+�~t��p��^��!2%%�%
�M�[�Ya��*�T��sGs�+	1�4�h�ϵ�A�I�Y�[���i�jF6D1����~�}�U��:"�JL���CMN-�j��3EB�:���b���*�����:���za�QzTrU��H����Z�ʀ��p��$�����[�١|�$��~���)+��4Z�>��P�G\��<���0N������I2����G�E�AW��6���������ί��=5�۲h��l��o���x��㉜���f�n:qLn�f�x=?�(�ݫy��sEE�*E��nM�!��q�l����:�zJ��7إU�S�Cx7ЩՌ{��ގ:�yQ$	�N���y��\i�J����R�"��im|����vL�.�I�x ���s���c���]��<&�\���G[ƪ�R10���p��x�éy��-'�d�̗�C|���-.l�̬�
f%�7v�����T��%T~"�i(Q��PjJ��ͽm�)�lv��i��߯޹5]o�$�s��gU�<r�cO>�%*w~瑣kJc{:J�}�����9Y���`y�lA4���Ow�T=�L΃N����Ǳ>oW-}�r�k&g�X�q�O=*xNG<m�N���NKn��'�����}}9�~1�,A�K�tt�3Ŗ
e��۩I��_�X��IMCK �byb��@�������`R��* _y�F����^�P/�F����e�f,d&V跛�èR�.��<�dX��
Nkg\��.��kwI�d�|D��U�^u�bd��mRu�\)Z	9��T�R;Z�
X4&�V��=�|0�Dt�-[0<ڪ=0�L��NS�T=�m�]l�Y���+J��M��:�A<�`rJbf�o`��@����Z��2{#�t�'�j��V�W'E�&h!j���,5��f�Uc˜ۂ���(iD���t����ݖ��T�r�a��-r���sr�SKK�]���$4s3Hs��f,2rs
��$�9���R���$��]��+��W�����F�n�ͺ����ml|��:y"�Md	��s�2��rI7ץT�5���dD��	��[cb��a� X8�h��S�Ĭ|gJ��%k{rd}b+B��C*o_B�is�W��d@��?Q]&��e�K_2�c(I.�e��C��,C�e�*	Mӗ]^ �è��~��϶b{	�h�Z��'��^�ĕ6Vs?7���M����kd���P�鉷�rMbxQ�"��o�ݕ�^Ei1W�c����L����8��t8�Y�T��� �\g^�!�A�}��umMҵ5%r�bz6	N��ŤL�(GBȨ��ܴ8��"Q�4�?��@I�1dӖHF�>p�1�+�-v��E��{�l��?�0]�^�UEzJ�(��Єi��3��8�ZbI�_?rT��s���6�+"��`.�4*��Vr�0�v;�>�ʂT%�׏7	�&�b����"��L
�Ռ$�����N(Y�[��1{��>�I
�\5��L�[�:�7�1%�,���)щg���G��sw`�#\Iv��g{g��&� �Ĳ"	EA���Jx~�Fn���xn%2�0�Ҹ T3�Vs��}|�]y9�y>j<���Z�g��l�Dț,/7���$M�n�&���7�q�����U�.�����	��z A����3Vt�z@���Q������>��.H�@Ek?u:�v�}��+tçx�ӏU�����qq=�#�)�?��[��Yi2���Ue�n9N�d`��}��LE���7
=�P����ք�,3Q��1�F� �WoL��u3mc�{)f�I���R��0���>Wz���R��2Gի��k婅��@,����.8��&M���S۽E�Z8{'�-'QM6j��.�7�R�� ���H��2E��4� �)1)�M�1��L��!�,s��[V$[�����l	9JJk����S�rQb���r�V�|k�\���13K�������
k�㓇	�@̛X�W�r��ȏX�k�d�l)Y���z ���ZxZs��_Jh�*�aj�%��t�gw'C/�gۢ���u\�B$F���2O��zagY����H�[ߴ|����Ji3�9%��J~Oʢ4����л֕�Oμ|�!�H��6u�av���u�J1�SM�:���4�Nhax-5�Vɋ�yO"\��X�d�QL "b�T[J$���C���
5�����(Gf����^�Tn7�Ze��H�(��)�M�dM܋�w�P�a��T�<+��4�Av{�H�|�9f�d�L���4]���'�$���EUM�9<N�:�0�@�k�����@������)���S�$K��LAӗbr����G�����5��t�'�̯LS�>���6�"�<�4Z��"��q!O��b��p���%�OD=>V;X�Ҟ�l����<ڈl�S�ۤ�U�;b�/����hJTc�A��R掺�@X~���q�p�|�h���i#{��%ޡ�g�E�V�&4������i����/"l��n�8ȱ��4���ٺ)*+L`�x�Bo����#IB8D�T��m,a�ׅ�u���x��M�CE�3�k"E�Dg���4m/Kƶpv��O"ʑSJ��Bl}q���ފ�O�i�j�����a"W|Ap��, ��˃��,�%WS�K� /����~s��.�.���!�_���Q��X�j��htǤT���aeئV����fq�҂Ct�+~
���o�T�W)o��L�V�43#im��F�&m9����҄W���>�U�]L�.`��cC���H���ШF�@6�Xs̏���q��x^��rW���_Q%��{���V�����>���Y�_�+!�qx�Bq�k�l���@z�fMک��#�Q���N���E$�:E���D<�W��2�Wֲ��C,b9���P�d��2�}���Kk�g/�����u���,�!��	����sR{��f�VJ�>o���MQ�f΢��l�
��Ӊ~J�Z��蛅�t�Sƻ"��'���,���Ua��H�k
ᒲQDf��j:���{@�����EA�히6pvq1����D�i��ŏ�wh�i,&W�~ק�g�XTCS�n��	4�(��B�A�a�{>��Y)�T�/B����8bB�K�,Q�ꆩ����y�]=zp����F����*qcm���/v��3����
�P����+jk9�  ��lw�N$�,V�d��{V4j]B%�(��=HMV�оZ ��88�7��al L|�r�[�0�%Ƹ0)�*0�P�>�Aƥn���o!��ܦdU�P PvX1܋�B
�M2�,�7h�:D9�ILt�3�W��O��� �!d�@G"�f	w���I�Th��>P��\��ۗy9䒥X�_h��ď/C;Z���e�~�e�W��<�t+e�f���r�Ɛ����|�ӔqΧ�����n���OzT�FT�+}#�S�Q�����)ߪ<��U�8�	��5�n|��BT��&����ՑG�$#$UG�Q�=�a��=�<u8��#��TqMn�?*`���Eu8�)y������ǒ���N��RJ�D)�%���1^K��H<#U�1<J"%G���H��h�����P˳w ���]� ��{��Ԕ���P�u�������ٽ�I� �!�ڃ\��O��XZ���>�[&�4����oO��;��žA˲����T��z�����Eҽ �h%��`Ŏ{����$ Y$�G����e0?=�n�������^������1H3�}X������;��s�l���c�Za,9Ŷnm����|�%��eSjߛ��������-�*S�Tl���D�#I�^�IE#&nq<��p�z��i'�+սb�P(��
�������7�l��D�0�o�lQ�����Vhx����Or��-�囯��k�y�Z�����%0�	���QFZ�F'�2�?��оTbya�s�ب(6^��ó-q}���7�h�da���>]>�X۝��獲�'-{����M�}��AG����7D����'���|%��v���5H�`�1����e�����ԭJ�*��ݝ��I�Ft�\���d�b�Y3�Ȅ��� #�u@;��xS!��|�S��{bi�6?nߎ�~���r�o@%�f���X�mR��o�G��"���S��R9�}s�����
���B��if7 ���4[� � m�
�`��`DV݆N��-���sô"��E�`,����%�k2�Uq��$�Ș�%R�|N�*8��{FD�&�>�O_���n����<��u��������W|�,RY�0}(�4��'�œ��N�u��J.�i�*���P8��n�\O�Ic��������|��2����G^��g�������+�0}��������]�I0��@�% J����Q�:�ڏYt��)��].�d�	��54�J1�#IJu�.�W�?#8��ٳ����C'�!9Dg�9x��%PO�{�l���`��,��zsp<��h�b�?	���펑�>��5_�6�����z�ڽoL�Kğ��%�y��㓳�3��^t�0N^�|�=����f�D4�F%����95��F�)���JM r&Ȇ:�>��R�*��r���� Y�b��7�@�����z��aOͳ#��@����F݊%��z=/4VmNOt5@��*��\zo�/}~k���_�ܩ<7T��Cb&@�/���+ꪑl��3v��W�}ϧ~���_8�=x:m�b�45u׏&/�\��,%x	�q+�rL�=~��|����0�ޫ�ˈ�g��f�t*7.�t�Chjg�&؋)e7?a�F�W��6Ǝ�՝��8���/���^��觕��A��Wr���6�k	?��������Ft�:��4πx�7�	�n8��͙ �inka���{{d�������<�cVO-�����|�����2�i�Q�XWe�9��ֿ���s�����K��Ts�A���_�a�u��H<��xe�ɴ`S6qQ5��,��O�8���O݋�����˄�������r?�}���������5(�/'����?���+&�d���m~Nҁ2Vs�bg�'BѬHi�������f�$�P,������aZ4��^Y�Px��Y%��]oL�2�������3H8���3���|��U}����9^p��+�f���9ņ��ˋ�ؠ��Dk�k')t<sp��J��d�cם�D��K�@?>�e`Ԙf��$U�~�K�͕_Xf���]S�؋>���������8�-q�M1e�������p�CX�y�|���x�l�\����� ��sp������\{x0�r^Xv�
�J�E�9���;�0F85Ӷ3<���y��$�S�D�Vlΐ<,�Ph�M�WF����~�w�K���o����w��*�5�q����:4`W��Tr�}h��iaak����I�z�,�Օ2�`�w	��#	���[�R�E���*��{�q��|����³4`U:�Z���B
��,�s�>��f��|���ZY*P��z�ӿ��a����>�-���KfG���F��㌈6�A����1>%��
).���o�S�nf�>%��Ǉ0{���z��X�Jzώ�E�1�R	���Z?[B�L�bɶ�~\K�h���[���g�
��� Z���Tي�����P���uWu����K��+D2,wi���Si�P�����L�
-��Aq���u����R9\T�?FzO��ū��c�CU������*6z"��9�[}14s�+�齱���p�l�gLL,��T�[�����03G��E$M�Ϫ��M�p1���Pe$bF#J�܇^��y��dJ��-�̥�iX��/�y����R�����w�Ig�Q^n&)��%Tl�'��E�"t���lX88F^v�#�HR���x��
���.�8!�{��?p�WW��uu2EABo9�=�k�DU2Q`���%r��mv&�ޡ��I��O'4�o��3��XL�2nf��/)�3��=�S�Qy,��Pyˮ5�$W��'��ʘ��a�Bra�%�b���*u	�%dI���05��U�AlpSc [��r�� P�����-hQ�gm�똡~� {�|ߤ$~̷�8q��&E
t���P߄;�(R�%��k�W��o���Z�Sb=S��Q8�e� �8UO��:	�P3gsA;eT�������[:���z��R����J��L��y�2t��L5 W��6*!+CKEiZ��0	-d�rd�Ti�>.F4z� yR�_���zt�L��G[�����!��h������������t2�q�w0�Ι�V1�Q��z|ytvtC�a;��c�W{�����d�3�pG��Cb5�
�"�2�`8"U1kR���x��'e�n�HPKX���4,�qo��M.�ϩ�T/%�Be������*r���wJ�{���_��Br[�_���`�P"$�����MIiH�9|#T,W�5�����$�Lf�:���Q��WWlbOMO�u ��p�<7���9�� �v��Pwd�ȖMJ"�Ș����f7���,U�"���.��lqyg��>�
��ĬB�D5���<�`�Ԥ��V�\9�-DK6��]ZKJ���j{�s���=V�=�h_�f`|<̢M�·؀�K�jq�sX�*���OÝQ�������f���8٤�.��+��X�VfF�o�������|�*Qhjʊ`s����i���ܦ
hh9p�a��u�����3��?�;����I4�m"U8����.������{���nu���	���ۚ��@1�e�Lc�6��%�	'$���\Sv�Ljۨ�Q�W�"x��H���bQ)%0�|g�+o
��&Ř��SVH��8���xI�������g���׀U.��d��pnY�wp��%��2�O����2
��܇#�����b�B�������o�>!��8b��%��_][�P��TǮ��c�_���,f��`55%��B���n��X��}~1R��Fe�xikѴ�O���I.3�<��	!^��_�Z4V�Ic,���>u��B��6Γ��Z=�	�`?��җ`�2wI~����u�w3��>�ٹ0��ߦ�{g�d����X�6df��Z�a��k�|�h��۴T���#�g�N]�������M�c����YTk[��Q�b;�|��Xc`栘�H�ޒ�j��m�`C(�'�͉����9���c�W���MȦ�k���H&fH�����C�$��_ϑ'j)�VX|��	�`Z��n:��o�[1�M�y�E�CEF�%��L���=Iv����H�s5��Ss�1Y�N�
[4�T�8�f�eӈ50Y5b����� �8�8��pa��x��L{�Z���Gf�yP�2UJk��f�\�=�tj�y�)%�˯-�ޯ��o\r�ՕSP8Y����[��K����Nꯒ0��d��, ���q��di=�%��6o	5�X�Q�m[�=�u�m����98/ #)��9�x��b�^?1No���%��L����µ����r��G�ڱm�N�Y?��3�R�N�c5��acc�9�k ���PĈ���(?��ֻҠ��"H��<U*8�2=�.����m�x�҈X5U�/�+&�����j�����l�7�.��gq�Pa�η �vh�"�N�uh3�qȠ����_ކ�̗��80$�W�ʁnZ!Eb���S��Ƙ3(x��D1�>{���c۔����7Hd��%>d�!ŷզY�֙�2��x�y>��L9ܙ�}Z�ʔ|�(�o��-v=�G|d���Ҫd3W����R����9�!^�j�U����|�e��D8WW����1Ս�j{�4c�ژ�'5�.yH�(|,,S;����Q:`��йw�ʩ���Q,Wgg�x��_�kQbR����)@�࿣�7Zpe����WeS,{u��ԍ��JA�&�n�R�cBF�yxx����kۻ�`�T�u׉ƌf�� �"�9�������C-�z���gږ�Ũ���ىC�	"���Q�|l�%5J��ɍc���tJN��xn"o>�����-����wybu�γQ����y���c:�a�B����/�)@.!�tE���L�l�'b^*n���r�h��D9�&v�b�y"�]���b>o�Sԩl5Q�9PZ)��h��ش	��B�rM��U��|�xMS�T�zqwshc�&F;&��(c`��LR��N  ��.5?7-J����ʗ�'�b�u��)<G�[F9782�����/P5��?M��F�����c~]f������j��d�����b�Z�������:7Y�;agb�jA��};>�9I�f����}qM
�,��H�sb��5͒�n�*��|���-a�%4
�q�vh��f2=�9�����[����u��y�1�����]���F�#���/ŧ����a4�Q2��b	"�/(�f�3d����=^���<�k���s��6TC�K�V��&����d9q�6��M���Y�6I��C��H{>�C'�x0�)�<�G7z���00��O��ä���CB����f���N��.���J5�e�U���^���XE�i�G7[�td�0�����u��1�0�-����W^cs.�N�1����@/7:�8;�$���rt�ŵ����|�vf��;��k,0�^�Q:m����ow��|���m�(�L���@��*�Ќ6��͑g�U[ұ[�����]ю�7�S�ä�א�Ź�u
�1���D�>C�pC���l�>��ʾ�{P������C���ڷ��4²�J� 4��d�y�g�Thlڜ�J��XL!��}�6�	�ኋ�5L�)`}߾�6��'�s���w�kfuۑ߂����	��b!�0(��*	���߀:��������%��o���AQ� �Z�7x}lttCgk�]��˓2C�m+M���x�bB?m�A����o��=��*�`����=��^HD�b͊E��?bsFM�c��F��/��YǗ}�<���y�l7^�f�=_[�S.SO}��s�i=��h���)FĻ@���:����W��\>F��Z�)�f�L(U6�HEJ���kֹ|ӳ�D�|��Y���w�T#$BF9��A�5������ � x�OȎʶ�͹�}�-��'�-3�,�|�|J��wU����k}W����E纒�	�v�w O�� h�`��q9"J���ᅌK����9�z~��n�g�Wz�������ܟ3.���t}���q���]�8����Qc���hj��p��g��x5�4M��r�M���MLPY��mn:Z�K��.��d&S	A�*(�}֎G{\�O��k�f��i\2�w�D�ak�W�Zy��?����A	�ߵ0J��`�~}Z���A��������p�z����:Rcl��{�wEx~X����j�2<x���9��>�q8�L�v��	/�s��eY�SC���;$k*�,�y�)'��N%<���-�M��"+bY�!)j�-�Q�;�|	x���5,
[^���'��������AV��Gn�z�P3Jc�S���֠�p��f����0b	p�+8� �}3����9�51�{E+�Iԥ4챼/؏>pi~Id�vXv��y�ds�{|V��Kߙ��o3[�3-� �_�w�p�Ϸψ�q�=�o��ui��<1�w���ik�:i�uT���,\|d�4q+�f���3Ԇ�Qr�Kw��o��%�qMZܵ��ɘ8�x4�!��dV+"�{��;wӾ=���i���m�C�&��5�F9��cׅ׻J�d������C�ٟ�����"�0ϕ�ܩ���s�����hJ��lK�1������+�k���=�P���I,��MԝEN'7�2�J����H�h��ֽۣW��?�q���
�5P� �{!�G�#�,�ש�wt�M����H��TϟVi�-�>drT\&hAɹ��؋���-��7�{j���u[e��lc��RL��E��72<A�taƸ_�����{'��=�����u�>�ݶ3��j>^��2eg����,���ysLxr"�hv�����FVi�d��ez�{{�'S"U�p���R*ɽ���n9�ݴ�1�iY��i��+E�4}B�S�L����Oi��^.pq����^���,��Ut_�S?��c��L�-6x�r��7.����pm��f��:t$��S�f�>��U��Qۢ�����2�����ǚ!�?T36��K?�v{��?n�~�q�9I]fĉ+{ݑ��=��#�� zPXb�2i��d�Xb�N9���3[�;��P���B�gGM)V�?"�p��4���Pj/5��oc��hn����9c��Y�k�T��n�4/���/��$.D��8f(̱��)u������@���l��M�G��������F�[t�_�COJA.A��1#�[�	���@�N����l���$��P��~� 7C�V��Tb!X�u��i}��,4.vʗ!p7(�K�X��Uas�Z���K��o� 7����͵�-��q�Ӿx�����Φ)���]�]#?�?-�<����r<� z/������c���e��w`�Ϡ13cһ2���t�ô� �[��q�L��t^��q�Z�6������8�e$E߇Q1«��U4�*��&�������vVb~�����C�������J����ô��ȿ0ĕ���ũ�I8�e.cF[�ۉ�l<L�/��h%�W����H�Z�?Rm��Z>,�|ǋ߶&��#�g����T��w��Z�?�����O�On:a=��c��\(a]X�F�!�6�ab���nzؙ�Y������SУ��'���dԄ<>�I�%��G]��Z��k\����f;��K�ѥN��ɍOLTqi�CxQ�FSO ���k�ʻ�C��'��6)o�2:�åF��͑Y��3���I��#��B����w�S��'ۨ�diT%D��'����2'!��?��m��yF�%uv�d�u�0�)�T:��5`�G�+��ބ�`�^�2�e;N����n��mh��;�Ȣ�Ӷ�(7��v}��{fYb&���#�.k>ETXY� �<�t�"^d�	L>��/3�w^W��pF\����9TE�Y5xp���%y
ٮ��3�r��XZz�U�vsR�\R^�&MKO/�_ظ��VV6Z�$ظ�,c��B����V��-ʩ�4�O�| H�\�)�3�� ������DδY�زs(�ӥ�D������~�;.���S>���e??=.���'t�rd��>6!G�
�*�d1z�]RE�jK���[�}d9���3Ȭ��k���xQ!V4Q.DV��ro���9���?��������Fz��?����"���P�Ќ���b�#��H^9I`�TN�yO�F3|��Y.V^e[[��F��VW��&�� �9�&G+Ǘ�x|�^��&G7T�\U��五�>]�^��8m�m��4��n�&�DBN1*^B��0�ff&g�4ҭ�i:kG��Z<0�z�I��\��O� t�F�Ф����@�l-���~k��.�Wd,ll��4��׭���!���ݬ`e �Zm�e�l~]���9&���Oz1��b��UӦ�1Bf�Zfi��"�1"��VR��c+�O
#l�MB�뇿�%����ã�C�?l�eP]M�4����	������������!xpwwww�|�������S�kfM��^=����?�W𽳋7�V�ީ�^N���-lŷ?��G�\)Av>D�umt��^����l'T}N���PIq� �K�~U�� �s Zs²�� gۉ�}�a�<��|e�Њt���5IQ�1�mk�Ws ���&�H��(p.y��p_�>M�-]�����
EMǋU(�Mhj�M�3N��5�<f�)��u��ʹ��u�	�<^��(������^{GW׬���t�dE��{|��f�NM�q��-�!��,�+�9u���T���?���0&lL�0���)j+ 
�YQ���b骕�qs�(���P�w "�OU���d�����#c:BS�/@��g�xn���"���\����ʪ`��瀢���xN�+��ï�sdI Zw�k%�؃2�PG
�^�P��Tŭ�諌{2f;nt�.$T_�@��[쐑��7J"2��1���q����U��'���d"��CaE{��h��kZ�z�z�>��#y�����PϩB� "Lٯ88���,
�v���K+	z#��0�rm���ˍ[���_k�0��u�Q �j���I���mĭ�K��BXs����+谑uh�%ɖ��W�������}��r@��+v�	x���-�����7f��gM�$B�Z.Ŋڳ�j9V���1��ʨo��F;Ѯ��m�?ɷ�_���w[�뿀M���:7��f�3��vc�<G?���~w=5�N�\J���̦�j8�pb{���h?E��Y ��I��zΔa9����#ĭ�qg'�9B�~]'&(@��@��A˺�+t__7����0�&�فP� ���?��%��;�[I�!�W&x<���(��#`a����q���c9�,�!��Rv��
�c�LY��-(ɋ�w�vq9m�rS���mP^9#'�h͈�r����"�%��_��oI���6��,QI#OiK	<�^u���vQ�>���H�.=�dfpfB�j�uL�E86>���T��)�F:�vI�Z��|ߝ��	�9C�ъ���<0~o�ϋ��e�V3�����v��n�M0>w<S�>W�g��;�����T�DEF_5k�9�(Ia�D����`�L83SBz�蛎�[[�v�JЕJ{�0�݇�UR�U������*W�v�G�:������Gֳ7����c�N�O+(h�L��>�>n2)k%�'p�g<�lkh�~�!������W�Ԝ�����L�:q����m�l�v>ޮ,L-�����?vP���B�Zy���L���_�</��o`�6�܅e�:��g�9�6�ҭN��S��p#k��d�
B$k�*f�Vh�R&��*��E�S�ӬV�$nʎ��f��,eK��y�B#�:v�qz��
ًk���1:���7��|[cl���j2Ԇ����_��5����B~;�[ɛo�'2����_�w����ȅ�Q\
[A{�4:WZ�߅���8M�̭h��QT����0�B����[��~���.
��~ED�mm���}A����T(�jmm�=�9�g�ON�B������FM��!&��2T�#��	���v)�<=)|�x�����X��%��Қ����?ݻ|�xҧ����<@`��P���76��x�[_��R�V�Ij�;CU_�
q�AЏO�d�����X�Q���L]yy�_��dM�:8,	�l���Vs� ���f^��k���|��9Τ�X�(|<*���u�K�U qK��3��9�$_�gJ��l�;Tm����y��&���R[ֻQ��?eּzQE)Z���xf�~W�Ss���-(��� `܄�|���<�
ϲ~��>��)�~���P�P]���3h÷���0�w�pQV⧦A��&΃�]Ż�.��kpLK��	�,���&��^.��نj�>�v�Xt�hL����w7�ve]Z�Ԡ����_}�e�+Ȫ���ɪ���o`NJ�SN�θ���ڙbG� �W�0��Ql�H�`y|�\��>�?�vuW7O��.(а�:�'�lQYT�{b���Y��o7a��Ru��EZ��D9����gǍ����ɹk��yDو�z�qz�Ϧ/7�;�Ztx.��`�V�E����NX&�(���!��+�lٶ��^J����G錸��K�"FD NπgЛa_���2�׿�YEH��h�2�[�S/ʠ��B���4f-�4�;<�[H���u/`����]�3@~<�*0�/��l�SQkvz�E�M^�1:�I���I����TK����q�G1�C���3�j��-r�\8���I�^�v�t���aj���6�sd�\�+�t�]�{�_���nP��}��}Mr���mx��^N��K:z*6�8���e���g��3g��m��JS@Q
r�sdC�b�m�@��k:udCc6�ED��׌&y���d[�mB�6�d۹h?g8y��(ʞ�uߗUhA.��i�@��/��Kss}���€��7A7�5w��r��#����}n���磷���	�3�K�.Ol�`��t�z_���@����$
\��˺��i����]|!��_K�EL58�h.���d"w)��9� ���%��-�Rԫ�&��3��~��°���R*�R��I�
=�%Ksl���}���R����i��̒���]�3���)��)�M�͈W�7�o�?hTס2�(gcp�$vgf��L����g\>jf}5B�s,�n�{{yb�-�>�"3� �0~����5�P
C��d���7I�	����<^Rn9�:gq��:9T��(Ʃ�aj�7�����af:��~ ���+( "�1�h�R�m=��e�+��]���~m��\�ř�A��ǆ���0����[��������Dz���ŧΰ�I�˷��p����֨��Y�?��/��@*�u"��w2i��ްlkZAi�*c���J��]�8�uv�H���(�op7�+��7F(�@_��0o��Yb��&Zf�=��a�p�SR������w��}�ز��������ea�5Ɲ"�'�hH�L�1�䂞 �����||/��W}2���E�[�)������U�[��?��\����k��F9���oz^z��6��V�2J���k�ū��Z��	Or_ٞ��\���_yry7���@�� 2�p��ٷf�����M��.��;I3�OOφWp��b�����t�Ύi�+#DG�lB�.��>#�,��!����3xs�'R����6���35�˄9�Ä��T���o�=�������uk]��ET+\�,0��ѹ�Kj|���6�k�^��j�uBu=	�[?��o as�i���qI�Vm����������sV�Q�mf�-����lp�^�z��\H`T
�C���^r��.��Waͽ�ǹ�u����P������m#��2�����%WOl�Wm׬{.�K�F0��hrsC|
5�fy/��X�H�����Ρ3<SWl
�y��|��Օ���)�e�¾�Ɵ��N]���r\.t�W�U�L����
w4�5�S����BN��``BCo�m��\��j�D�_Dl�f!���~�� �Ib��'eR0J$�%BY��Ԃ'���(`�ӹ�"�Ш�gfwG�4:(����&\6���	�/��,����<�F���DS�=ꏳvc��g7QE���g�a�\E����?���$s߱�܎�͟����=6&�:�<����n��
Ɲ�iJ�>�f�}���j���y��"�CE�m�0f( 	>o���cЫ�iƪ)�e�m�Д��EH��=}��	c�e��^|�K��~sK���v�K(����n>*�4/�>�`�����EBw�D�c�ch$-@)�g�Mr�!e�_Ǳn���"WZ��w2�}x~�!�i�Ƥ��p-o�}��v?�9������Ǜ�3ऎ�<Rl��p�x�o�O6�~ȗ��h�w<���KO~>=��>�l�:]X���q�7�dw;����5<�^�O5�(W��C�B�����4c&6kY�^_)nb����,ϗ�3?�����ڠ���bn֗����&)��+��zfјl�ݲ7���SF���>�;zG�]Ɂ^o����́���/#B?]&;^i�>wS��ڠy',��w�D{LO[��/�/Wl~���ڴ��g=�������h%m��ǃ��H:�GD)Ք�#�cc��ޅi�ʾ����)�f}�.�J>���{p�~��̇?��>�Z}���/d���CCx�Pz�d�M�c��g2���8�,�|ALh�_z���a�4�U�Pо��w���1';/i-v,�>������� �Թ�gm�kpɺ1l[7Y@��������T���I�w������G!���a�ø����#�'��s3NqER�l�C*i�A3G���N?O&v3��_����՚��CIY���L1�y\	�@�󋢖�􋩮n]焦Vޯ�h/-Pڥ��6^�	vs��=Δч�3!���j�rP}D��J��I�� N�f���H��)�~Wv�1�J)���M��V�燠.��I1ɿϧ��Z�!�%�(�b�����7�v�/R�)l����l5>Ā�_9v�sw4��P�N�{_d��}$��U�it,aK�(Ֆ~��դ�����~+Yͺ���i��L'/=ꅅsҕn��Vo���%G)�q֏��
�BJX�ُ�P�QR���.>��چΖT��݁��X�ɔ �yh��ZgtS�zٷl4��I�SPʠD�/�	�Tc6^��cfx��G���6����f�_"���5���4��A� ��:y��-Z�R������'ᗐ�h~DO��H�i-�;�%�L��Z�����|��?���d"���X}Xq�rf�*��4�C~-Qߊ���e)���ˡu'�RD?<��C�<�i��^*�=�x'k1 �Z�1��*Ü~G�[OM�y�m�_�po9{��L��_<?����P�'�ꔆ��Eq�[j��#�Z�߂�!-��㈓[��K�{��AY��`g����6DWyrD]�-�N�N�PޗM��V�^=�Huw��u�E�*���c:`�:B^�jr_}���C�2d���� ����ji��͐#��J�����QY�X��22"�����(բe��ޑ�͊�Y��-������f�-�!�x��6�;�֚��"��k�������Mon��M4��&j4�����p5 ;2NFܲZ��H�\4�?w���N�Y�_
r ���@7ő�z��}(��F&��5+�Qi�8� �1� ���݈�B�D��:��h��@r�ۘ\Xg�	{5Vvǎ�Ը�_�]��1چ-ԯ>�g�Kpa/ �u�c���O�$6C�_"ɭ@G��d�(����`�{�W���]�iҲ�y$�`��3Mw�w�Bo�ٚ�c�ۗ�?�ient�`�-��l�;eD�M4���,  ���F�\6���6�A?H9heoY���n�,;��L����B�OeaV�o��Z�n�bu2X��t�<Gbd�&��ATbͣ"�ʢ�H��2���Q��Y��K�y`:��~9 ��-���׫$�C�X���PKo��Θ�y���,Ȅ|y�M+S�y���?���,�d u�U�N�5�����'���V�8 ���Ͷ�*�/}V�K�)(��\���V}k2r(���t	�� jZ����3'�tRey,
��"K ���b
i�c6�_��P�Q�S�!�ٞʕ��q��~������Y,/���"an�挰񃓱���fcd@�߉;�tE'���5qG6A]���3h3 3(I9d�1=;�{}����k�h�J��� ��[V���1#�t����:Ǿ�5�Sequ)����t��NR_QUT���ravfs�x�0
�!*QXD�i�M0DT;��ۧ�r�*�w@Ϟ+>���B�[�;���~@�C�q`����aG�U�af����p'�Y�i9����6YCW�\���W�0˫FOB����k�+�<N��44�q����E|[��žke�ԙ_�:��;�Bh����7kv��qgqmh�H3�{+W���`��R;N��3��o\3�Q&k�%���;Ȟ�NK��>�$�pZ���n6���+(���{d{������?��2�;�Æ$�j�1_��&��O��C�d>�ujGLSM�j*ݬQ�8��Y�9��V[�V�XA[{%E��C��7a�qʣ��{w���` �*_+>~ʃC��:�R�3����p�ם:s���
���� Lx�_;y�Z��_0w����!��iD2�^��g��Sɔ�qA�o`�Յ|��X;���+�*wq�����FR����j�����V��R]�6&�#{�<H'�Q�]T�+?H=Ρ�z��%P��EE�2�%VeL(l=���/@��V���s.�?Rb?��&C[���%��sw�C)�e�������NR�+::�|�6H�^����'�U*i�R��g��i�EAabzq��l4/�/����[J
��R�c�p���8����k���� Q������8�^�5�z�����`�Kx��"n'�sZFN\|wΟ'U�o TFy@z�;��Irq˭t�m��E=�}5�� �(�*T�hqe�(MRx84�P<��~�dqzH a�|?�\o�!�MM�׀��jt��~��9��m3
N�AJ�H�!�(�h�j����u!��:����Ry�J�V�(lq�#5@��nB�My��'B(��:��)�Kl�/x��f���Q��!aaMM����3N�zu���ɱ�Սu��w��K�qL�𹿔�E�~p����dnf������o�-�X���w���.f���j~���:=���n��.f0Xcw�ÛI�@�Z@q<���.q|\aQ�fi =M^F�8�����p8	�O�b�m�͉���3������p`�`���(S�d���d�������MfU[97k�!�/Rʣ@!ա������R���f�4������z�=��'�w=u�`�̉�0Re�BBD�seO�D�D�ʈ�g�Lb�_2�b���4)k���C֖c��-!�����E�>�uS�mT��O����w�S�V��>J�:9��([5�²���q¤�>�ag'���!��Y&�o���-b@>9�y�F>+�w�FzA��
��=������'�M��)dcgg��#<����}`�'P�&? �����ysr��H��7����,)�D��u%���,^�"��j .���]GP���ܔ}��
הM)`ǀ>�H��� e�S��b
c]3<���|hHyV�7E���r�0�ה�R�@��F���UD�ʟ��3�	��ϴ� ����K�����f!����Q
+9&��|�3䰑��4Bdwz	�W7C\^2��g%j&���TL�c؁J�{Ϣ�%Om�T�H�?Ū�$��ʴ��gf4���a�UUA>-�Δc�Y��E�}���_ �c��fi(�@7i��8�YVJ	S������Q��4k��~%���M\�Dd�	y�������J��KG�	"�8K
���J�=�b�=No��i�0dG*��j�b��\��iz91=�4�an�8K�|F��ٵ�d;X���,-݀M�)yXz*�Br��8^�N!'�(��Rt\���Px*��N�e��'�:�z f�͖��<�rh��(��k��⢍�j�7��z����g1ϫK�[W����0`���/�?�-��l{?Q�Z�.۞q]y&�X�B��g�A:ը�	�
��u�$����$(���R���`4Ɛ��ʤ5z48�������y�9�lvy=)����f�ަvmO��a=���<��Hʚ��	�H���|d_}1�-�)��Dw#�؞3�:0X�"k^�R�\ā*]����M��r�
�G��B�prpH�= �Y�bmE���9m���d�ഺ�06&�^X`���9�Cfn��F~?�k+/�r�͜�)�~�F�GD��}l+�U�~[��F��tԙ�
L�2p%�9�+C7��4�F%�^m0�<�ȃ��b�w���K�Ф�_of�6�twW�}���zDҖ[Q-+�a��X�Ex�s��au�^L���_�x!3�|q����:G9��]��FO! �*\�J�Mdzc,�	Q����J�bz���@4���o�I��N�u�k�e���^�������K:l���m}	M�}FО9�[�I����\n���9�����x���ʟ,j�Mx2���+g9�@��{#OҘ�W��d%��cG��8��R́@�}:�,,,SS��iU�R�`�p��%�8<a����T(D+��ə�3���+������؆��
1��U�5�+��Gl�67�X�GjI|'kΡT0�� ��Ѕ)n�v�Y�!�\"�R|L���(�lx���'�J9%�F�-�}KB���=��3������9؏?&�*7�77cy�* �\-��RUb��n��Q�Vӡ/j�/�[��m4_}D!jxj����Rƶ[��w	Uj��_���ɑx�r��HZ���OR1�U*�X�B���6�{v���7#I���'Yk�گ0x'��ur�������ܯ����ó<��&!(k��=�Y��F��L�����A�6"���8!Yc�0�2��%Gkz7�菦�2��ؙ������N�y$��yhqd�@�2����t�c�]��d���7@��d�q�%�3��)�0ǖ)�c���Wn�����y3�63��Țs���%8i��5���#������@����O���oj	��Wب.��@���@�vc-b4�I�9�/�XS� ��ѐ�\��O���]p�������VQWY�A�����`��n볯�nMX�M���>K��NS�A�*�#b@*�?%�)ֽ���I��y�m7��X\�$#^�	��!=}xM+K�\~��&�WU���+��-<���ѺjP�\�ͤ��5�馌q�X�I�J�=A4	t&�}^�S�I/ԡ��2{GprӍ��&!ֶ�,�o�����S;b�>P�����E(ݑo��|sU�ӫɸ��7��߉vX�������x���M�Q���P=�~t%��f��a�����H�f.�a^j�uF�漜�c�;:xp�!x�
d�#�w[��y[��l<!%�6TײW���e�ߑj ���<6��,�4��G��B��|��]`lT��9D�}m����@�3�%0,�Վ��:���Z1��P��.�]��bj���V>ǲ�̘�����L+-����<g��&��%��:4܂��=��?�}���h5Ĕ,��nX�������vfN�Vc#�ޚ����� A^���yW\2��	�&��85G���_>	;�O�n��;#c4���F�j�2�rHJ.e$g���hc�2&n���6�_/6��}�,^�9���;��R�p�.�{B���ExG�5����B��;�Fo��/%И����fA��9��ґ��wb��.�5�0��id㮍�#�8E=R}�k���`��hj����Kv>��UesgL.�_���U��p0��h[��#z��}M[@�G��@T�v�c�[깷LbO.r�/���+t���;6%�ӹ�4��i�_�ZD��9	`�B�^S=>z�����k����M�~V�"��s�)��ʋc�pi%EC�ϛ����ʮ�m������(<�� ١������g��(�X��b����t�R<|����n�ֵ[0��0�~�6	����1�	f�m�q
yo7g9�i�k|�K��,29�d����b`B?�{����`�=^}�c�Ң'&	� �S��{��*L$;��ք����CC���	x"�/[�B�9��қ��IQ�i��bdP=�ZY!�J�I�:?'N������_Ǘ	��?r�T��>.G+V���6�� �C.A��i�^�I�Ac�Uj��A�>ٱ��A� x�%��
a.�D�O�H7)������z�p�Wj�"CI�����y���1���\:Щ��"���[m�7�(Pʈ���e9���-�!E0�2�by3$s�	���߽�8��d�~6����N�2K3;@���
��H��1�����C�B�rM��blh��� �A���@V���Y"����ѻ�f��dI�)�QRn#�a�t��J�{f����	���C�곈�㖈%ѩL��	�U�P���g�����p��嗔H��a�i�7{$ȔH��7ܻ����x�EG��c�E�x�*�I�P�(��|E�#���m�,�#>̅�Å��*W��>u�ւ���HN��Ԟ� 7��B� �RżtL������K�g������.��VB���v����ڄm|� OC�R���v��c��`qU�F��"�p3
�j��%E]���XX��-�݆R$�dr@Q���4#�-�=�& =~�)�#�p��e��e� ^�،��9�h�n��~�rQ���&	n */�ݬ���gD�f�4�Z����(:�Nh�y/��]�ػz�T�x�#�?�։��B�)=���u�eт	��*rPfS�����O��W�JӐ}n���d�}�
_Z�5f��}F�Kh���ri1�#�a�'���rO���i\�fo?y%j�P��1�Ou���0��,�mMc�z�r:��蓜q�A�����.u�~^4�b.��. m����V����_t��4�饌��o`j�g���H��Ɍ^ZQ��%���0���iϒcN�]�i���+�\��-�xu�:4,�SS(} r�P%��8&������f�������hY�e��~�5F�����Z�5s���!���E���)f`[���7��_\$oaG�K7����+	���a��(%����7�ׄ�vo5�ds�>2�ӻV�k�'����cǽ��}�?djp�v[����w�(�o� v���1�oh���)�z�����*�- {e�=����o�d�}�0�y%d��LP��"�W|�1�w��c���p�M��������aW�L/%:O!�F��F5�;�*$;mE�+�A@/��'G��ȷ�`̎�k��ӷ��0���E��|a��c;�}��bFKj��������U��_=���G쫨$�yxC�'X�X@�ճAX�2���!�K�r��jŕk���t*��J��v!@����$����Eh������J#�#��s� Ӌ���tC�q2QHj�i��r�D���#ʖt|)�$�`[lLD�������EBȟ��4F%�<���P�ؽqJ�0{؛C��1QiO-�V0t�,C:j=�V{б-wm�/��60`���O�m���#��^D�{s�ǻCgapS�	}5�	���x�li�eJaY��G9d��[s�6�d]����@����+�AR�E5��(Y})�k�ڪ�=� '�[Z_��KS�"��:9_\H_lZ	Z���N����3I�t�đf����C�e�aa��ɼ�+�LQ�" �D��pؽ8?O�w��H�I��؍�t[|8����� �Ô��'UF��I�ٙai�4\<yY�"��ܥ��+�a	�
Bv�!�����]@\m�u-�R7S7Z$������H(9�u} �1���Y��k6F�Z:3p�Oo��(d���5p8p�}��1}��rtU���ߦN�'?�VK>CP���6�l]��)�b��꽥zb-�0{��idx9bjqaR�x��
����"oq�.�Tn�/Ϧ4@����d>����r��[v���T!P�R#V���&`��ʤ#Vϟ��*��\�X8��#-�r�)�"*g�ݲBNսe����f�KISQ+ý�������X��wP��M�,�,
[����c��s3�2$F�N1�ZwX��zzug���lW*mS�6�TL+��[Ȣ��ґS��v�����W� ZB�xs�Х +���@�r���#=�|�jHcOf�@?9%5]�5d�{��U��-�ts]�Fm�o�u�o����t���k����1;N�*�	Y\�%�MGy�f�:m�5c")f�2�I���孨�u#����d�1�s
.�|��N&9iW�N^ȫ��H'�gP�w�_Ӵ2��.����p��+�oH�&�����\t��5)';>�ds].����J�"�4|~|�:ғ#���E/���4ؠ:؊Ƃĺ�t�*�a5��\$�X�&E��|~����#lS_��ŧ$�(�Ç����t(tNQzA1�\in�uAZVJ��!��U���m���I�_��Y3� ��u?�Ќ��fn r�K���)�z�C*�p�̢�W���ڡ�NcN�	��"f�I�x/�(ϛ��#~kVJc����<�H(��p5��v��R�VN�h�eF���6����2E�dh�RR�O�Y*�\�@�H�S��E���
�UH��ז��<��,���1(~G�T'�T�����/A����#���3}��.�=Y.�#;����[�b֡�����l��m���t��:�QձmI�X�t��� ���+4�!S�s;@�άؼx+�Ҡ9�5���㔫+~cr���YB�{�DE���w���k��q�>�w����;��N��}�g1��"����L����<��0�fN�ίH��_������:��wtUP�"����'�[E���9�Y��в���uc���rd��)p��������]+��RR��������:�5�J�?"����M�1ܢ��f;�l�֥(5�G$?�g��P8���`hiy���U�hphU_�k1�>�WfGv{���`f4�\�\��
�:�E�/��rU�����eQX�ڼΌ��"�>���^�*����J����	���8eͣ�9�+�f'��U$ UW�/L�<�R\ٍ0���1O�W�0'h:oTQbn����;�%�q9d��]o��ZƘ��|BSwkۍT�����@�l*�	�\0��������:��O6ߦo�8�+�̐����͙�N3r--J/��qw.;gb�b�o�J�CG}����*�lC�t��MA�u!B�"�N���^�pSƪ�_����v�a�������ߡ�B8���#����Sb��B��>;Y{��l�O3\������� y�=���v�4���?2TWV�b��Q4@��&�ҋ��k�������S/�v(�{�n�Փm�u��r�/5����wԵ'0=�@�}ٖv����wO[
/��.�?I�ߛY�7	�L���uH���f�}Ip����2�2��zt�g��V���V��I�Ƿ�~3��͝@��6Q~B2$����Z��������|���;P��G|��>ʨH��.�P��xT�a�]}3�dL�ѿ���xI����O��Q����CRe{p�:�I:t$��?��{~k�G�&(/�6c��t��K-)È:��zX*���W�o�
i:�7�ћ�����ջ*��[1ؓ���|���:��>:��54D�?��3-�n@"ۗOI߄�S�RT�ʅ9P��*�R�YC{Mb�h���c��Q:�|BH�y��+e����� �8J|�&���m�~
��2�F�G]���7��3�}RP���q�"H��|��������uv�f_DI���^�Q:�;T����$�gv�Ǖ�n[�����b��2q�����1֑^c��&!hn���km�4��t�'� {��W2��3+ǝ���+�W�ٓ-Z�`B'�w���ߜ�X�%M�Y'�n��!׆�:��G�f�v�ߨ�I���EE���Gp9h%��wn��P���)�����%��\����*mCε��8�w�?�P�0���� ��
6x�c��fn���G�|�r�r���_$-Ѣ��*����k�jwc�������E��+��7�ʭ}�*����eR��&�q@-���{��d⟥%�_!��s����ݢ�i��*(n�S��������6yN@3��Q�<-��ؗ|^q�/��է�z'�-:�&��.q���l9���_����=��b��bG�s^����^��	B��z=T�yl�����~��<��b��/�_�
:,���K��M ��j�z~��ޗ@o��~�s��:���תM��g�>��c�	J��`�=I�?�|B��dddY/9.�B�3��t�@$A�����8�a�;���͹��N�V{�ۢ�vk��S3���B�3���Jf:x��ݦ�3%!M\�d��q�_W�= ��@d�d2���
n��Z�d�eΠCkR[�>�ne�b�6���u���_�6��O\�z�G�h5̆�<S�ͽy����� ��y<�X��庡����Y�l�w�R$k�*ⵐ)����;�:F�t���T�%!I5�wgT|���Q�u�����"��S�e��^�"���Ne�.R L��1D���VKq"������L��$��Jk����ٯ��$d̾=F/�<�ˑ��_�%L��5VRs�~��`�R0%E��<���*q�_$Y&܁:F��*�҆/2T�����/!;g/}u�g��:�9E�k+��L������MEZ՜%����+Z�������ft�.Õ�+�ͼ�� �V=���������d>O.�35oe.��"�Z�#tp�؋��t�/W�{Z-��v�����q�{�@_��#�P��)q!L��_|
a��N2&��>~����~���o+V�^�N@d���Ɠ��2�y�܈(ފ^$8E��01육���<����S�ʏ�%��լw�NG����̐������P�ǐ�~���~�#x��4������<OP���t�~�r��~���)Em츪�9����`�4�j�r�X�;�T�=8��&"8�.�Arz�S�y�B�P"'[1�O�85��1��o���)H�E�Q�X���V�:���֚�}Wc�^U�/�7D�G73���:�#P��o^��>1x�>+�wH	�Û�+לr��
�r�P��+V��}��EF�y��8-]N�B�^f/��_A{�&���mCt�U%�>�5�[�������k�D�Q^ʭ�r�O�<ai��\:����]
�w;\�����-��U�E������j
P��zO�{�\��$f04.�����d])x�4�Bc�E#��������
�*wH�"�7M/�5�"��NN8�s���������5MBoo�y]�߄�.Rz�5@���B���0��+��]s���>���'�4�VꮾT����3��p@`�t���r��^�X �Dy\�9�ov�
���8\��\5+''%����z~A�۷$�e���0�<)s{B������MaN�+xV�T������8���s�����1tE�!	��m�1!-�����a����C y�<�"�$%��$�GVVY�|�29r��
ZS�ӳ���ޫ�<>$X���a7i�i���f�������r�� �r�6�1���yD�-}�W�@�>�'�O�QV�eNpc��Y2g�џA�4ƌtf�ġW&�[rDK�K�[u}����Y�M�&I�1�z�u������ =�b�/�76v���c��=HU���V�b���(���"�V�3�u@ʾ"��e�u�l2�*���K�a$3J4�	����?�`#d�,�����'�gj�	��*D���?~˫�	פvԛ����F�� �/P�#�
Z͔�r�E��-it��G��IB���Ǻ�xU±A	w¥t��rl}�������B�^�,�:͍�q!���̧� {F �*K�*ƨ�x����򸰹� ���_�}7��^�I �~s�?�ۺ9�	?q��f�?�,$�v"W��B��r�2I�2?c+�KZ��Ʒ��RDH�������0d��\yon�ŒV�߭b~l�����T���	[�h����FE��e����-"c�	yp���I�𵚰�qN�bvЗ$`��d謍0b������0�P��8*�
��*4�h����]'���Z�Wo����s��2s�?n��}���>����#�Խ��+�
��j7��Z0L��-���Q��7� rF�|���+�˥� � k �P�P,�}��׻J&O)��܂3l_I�FbJ`�#O9/��P�Q��a�L���M�j��޼���6Q��h�gϯE��O��7�D �'3��n��lY�>K��b���BkUnܞ�'�w�<]���}=6���
�f�n��[A�,
h��,�k�--��5r7����Qhi}u��<���Z{f�y�L& fR�T�0q���]����SX�7Է~Ξ'��Zd�1��1g�\��!���i^L�:S����Z=��]���>_3F�@{fCv�v�G@\V��,.++��E���#6vz=����OHR��)8"`Z��J��m��5��#&Xa�2�QAn&Y?�!�*ʧdw������:��,6i����nu8���{Ֆ�m�t�[�����:ٮe�n�:�Ʋ]�g���=�}_/_K��\��;��'�7��Y�hVhDy�}\.�(�]�tT��q�|��$�������-��~��DIƬL��+>=��/j9�r�DC���[e��$�ⷶp���.��'��.���aLDٌ?hLL�W1J��"���߿[�H���UWu$��9�h����:�"�����m����}�6J��O�2�2���ۊ<1"`V\�3.r�18T0[Z
���.7�/�~V�B\\
��-�T���5��N+?2=z�؅�%Em�iG��i]w�"��O �KI����z���V�*3}k����;���b����d�g��Z�8�<��W��:oV���,R_���~g����>Jc|�-�"��U�/�Yw�g}w�'�z�nk��u;fS�Bq��j1��S�����o(�]b���8x7�1i˹�3����;����.��f(`'��%H�yFx$COLr�m�?��4[� ܻJ��zi-2�G�{YC��hq̌褛~��{���3b���=<�`��Z�X�
6uHJh��$��ϊ�:��M�
�@n��J�|�ZF>N$�ߠ���֩�W�����߹���\Ϣ���U��ᭋ��"������(���^ʏl%�HD���(�P��J;�<�����~�7] ��Um��zwG��X'u(SyGLV����j��^H��T�vߝ�j%}{�V�ld9����	�)A&�8M��S�<o[[|����羜0��ƁB�"�Vp��ˡz�!}�U��cG�f0TX�bbG�_����X��$62���%��`�5��K�:�aҨ���5�Vh�8�hJ}� ����p����ee��U���517
Un���P�<.���"8��8��eutTJO�iR����0��K\�(�8&����Wc���"S�j��rs�z�ֵ��>A�_�Ȭ8K=�$$�NN��E�¹g��� .0�FUd^�<}Q=��ej0�)�W�v��[
oySMUgG=^�Jz}U�Fـ�v�aN%$�P�_����_!����_����H�{��+��E`I~�|���t�?	1�g�'�����<D�겾+�	7a.�=���0��D�NI�ڱ�,��gI�����C,'NA37�G�����P��le�� ΃_Ϝl����(R_H�c52��X��(��>ǉw"���[o�
܋�H��t
.�)
���Z�LU��ˤ}}yyM�D�U��]�X���o>�Y���9�6�RTD�U�.t���Ii�}�yQ]>ś+��5���H�(���h���?z��4VcmwW=q���p�P�� #'~s��<����[����W{�v�啓������;��ϡ�k.�N�R�4xH�K��X!�Csݸ�!�WR!����Ȏ�,L�TptX)W�i`�b����_�{���(������_r��[�{M��qe�J)�Q�7��[�E����cE��P B'	h=g�'��~t� �����8F�����n��3U��Q,H���&�E��v����8�u`��ִ��`�:��U��ڧ�-Um0$X�����[��E�h���u�R�d�(ʣ<���]�m��6i���ῄ��a�yS�&x�4��y&�pc����'fi�4�f#��88~(j�z���e5�b��J�ά�Q@����־�h�$'�V�XHC;[�Y�����}A����Rĸ����%�P���A�Ya�k�4Q���
I��o�kd�df���LN�Z?#��5�M;N��B6��s�O&�-e��r��`%>����ؑ�Ƽ���fܼ��y�^���� kmPI�	7ߵ"h��Ryh-(i��Z�O�;D���C�Hb�K��!\iĄ� `RL�g�A�5�;(~�pw���	U/n}�&y�]��4�$n���ۖ<�Z�8.���Π%ږGS��!{E'�J�o��V�	
����GN�DHFK����z�b5q2eh2J�d�M@��,r�H�v�HqA��x�� M�=򤨫#��q�J��gqݎ���6�U>>1gV�~фH	��+7����u�80M�s
%X��}B^!Qn��K���r!����U�U� ��̫[�")�IE�/�m�v�:�?���+V����=LJ�DP@H���GD��4���H����c9�@�'8�1���1p����wZG�{��iEg3��
�
Sy�FdvR��w*$�T�K�VjM���͑?����.A�g\��C� ����8k���.�kC�â�߫A�������)§UUp����~��4W"�4�=��S�N���eL�*��Z���Y�FT�O*����	�Ƅ<2���F�i�+K���~��őTC�Ƞ�U"�M^��Ċ�}�C3�8j�;�n^M�U�]��Sx(N|�,�+9��/����}L�8�rw�N�@B���5uix�@r�:�>F{�R�d�B�7�l���Fr��}�y�X����_���0��
��:���ʹF��MCk�àN���1��]nM*�ɴϣ�Tp]9g�D�t��y�k"��z_ܽS�;;+�0�'��K^�OZ������O�xf,�t.-��Tj�_ꫭϲs�;�f����-�p��^Ƨ�� m�:[y>�pu�2��X�j�`�|G��"����ǌ����˔\'䦘p�A@��G���G�wZq�ʴ8Mb«$��[^HU7~�U:�<ʣ��	�9U4�]B�Z���%�3
�,�;��撛�w��^�������`��uD�y::�[iϮ���c�����q��|�w��&���^v������������Ę����'�^�(U�@�����
[�5�1ڽ�A	����[���>9�V&�.eF��6��4�����-�$A.VN���e��������{پ]��j7�����{��qsճ!/I�?�`Q�N���5������:C^�}���Ō�q�c�Be��o�����[���e녶�8_���;��o`s��6�4�=��ٛ��5Ez�RjV��P��PV��O��''�}���@B����4{���O6�A?߫�n�~�����8���Y�5VX�#������vu4��ZE�A��YhL٩f9��e�^a������=�D���:�����AJ����^Vv�>eFhВ����������+q9�����H��k��=��m�E� ��J{��ǉ�e_�t�+���֞��T��������ׇz�{�ZN��.����� Y+��щ	�l";��9j�����?y-rM?%ȍ�ͩY���_�<D�d������5f,��-[CE��C՝Y^�4�e�>���I�n��&\��
�Nہ�=��ӟ����Xǖ6w�o�VO˺P������I�Cq"+���AgP]I���G���������he�1�[:V��~��h��X])��z�7������]�U"�u'7�,��x��(�t��7�AE�kӰ���ػr���Pܛ���:O�ER���!�ocxX\�Jbu��u�m�?r2��w�/i������. NJ�p�ۑQ9���
�?���?릯z{��xFҏ�����:�.&s��-�!�!�,<�*S~�=�'����ǖ�fi(��-��C��l����;�d䳴��HG#�ٜ���~Jv����1Q�y��s�D�j�{O��!�FS;��%o}�I�Թ_��v��m��`�yW?�ݧ�ӗqo<�����W0n!���I?�XBɿ��EX\BSǳd9^���<�~ �O���!�i�vP�����fF_p�(��������~�z�S�������MRnn���P��%�ń+ ��4]%m��a��DG}��cףߛ'S�b��G<��&��F��>����֪ܿ
�=}6+8���E����Z�i�xŚe{3�c�D�V�d$12Д�I���RMF;�⼷7K�z|��Z�6���~w*(g+��]�/��aB��6\p�����}�Z�~�95(`��7��Y��r�f0�"�uܑ��F ���D�V�1�p�ҌB�"�93_�#T���.�S&º�rrF����_QE�4���=/��п�{�2��Pݕ�����^i�����~N�st��g}izT�?������_�*ف����b+/�e�����nߜ���7u� ҍ*���A�D�g�(��ˑ��[�k��U�Ģ���P���Ȧ@G�'�a���,v���W@�5�$�}GZ&��*X�����H�dx�7�����-x*����# ��<0O�0�d3��>����j���IS�A	���\���;A���M�x7��x
��u��|.ǷD�y�.��Et�b7�Ȧ��5/���K�n���_5�z��)+^_~�X�c���E�C����߲��(q�O�=��N�$2t�=�g���!��sN��N�`'�x��G^@̂��M��P>�XNC�T�ۯ&6|X�&U!&���-��V�S�v���qt��y�#���7R
�e�-�9m���L/�I��C6g�m��L�2�!�����ϑ���
�yk�Nb]� }��.j͑�έar�#WT�����S��\�����	����D5�	h�ޚ�7�F�e���������Xdp��ą��ur���-��r��Ru������<��&H�!��:��n�ˑ�ZY�~q��|9�p���uyw��2S�W3�)�w2��_N������Vt���̕++Ktq)J��������Nu�����m��&v�
��ĄR�j��R����tEdm�,���z��Xm�Gi���^�B?�U��۠kbi�w"���#�*�hҥ"�3^D>1��FﳂL������������@f,q(� 4@�g=�R>�6���ʹ�nT�OJ�?��w�3̥��|��'��%z��y����{���4j���������z��
Hf�L�����US4�	!(L9م=B�&I�I�����Y�l��i����1?�:���SN�u��������X�n�wxI�|����X���|�lY��ME���E
��h�H^��O��P�3�'ɀ�g'\(�����{����Fp�щ&0�y�@rr�q�5�S�S勜Ӑ�̌t1&�T�gq�d�x�MU��]f��v���Ȯ0T��+Zb �ݔ�G��+�8f|�X�
���@T~r%�s�Z!���Y���)�p�U>^S�ؓ�|qln[���k����l�T�����Z��m�J��;g�ܲ�; ��i�7�^������l��/B�h*�⁎��gNv���_XElQuc��N�z�;.˞��9"���D���ӳ�9N�.m7w��O����K���+s*�f�Q�~��v���m2��]mc�j���<3ڤR������֗E��Z�(�~�7���Av�c��,��#,#DN�8�|�d��2�r�ҔX)�=�τ��T�)�
�%�{I���8E�X�SM������*dz�K�ʫep��u��(N�J+Q.��5. /�*5�͋�:�䚳a���Z��6��H�z�" ��ڮ�a4Xi��nj�ے&�D��'ض���N?��ۭ�\#v��%mķI"�'?랚}�ķSK��b�O�!��'��'�
�S,	h�0�1��U4��!��bUo�,_~N-�LM�dāo]⌖��O��*��&B��6��)ҍ�K�O�ѓ/�54}��i���<D-!m���*.ϋ��PB�3�����V��Ĳ2x���L����<����� ) v�r;��l�ܷ�i�-�	�1ؠ��,v��!�t���^�'��^�~��-�|,�_Mh���f�s����vĚ���2���z$mC��د$D���m��^�<��Vt�B�А��8M	ER�:�?��7��,廿ki�;�IZ�A�kMt�5Ȣ*�A�{��)6� �w<��*���?!����>�3�yz3ab�+�=�:�(9�(C���z���Z��Ȑ G�����s6�tg��B����sbbZ������WH�
r��y�jE1�ܔ񦻭WB��,��ˎR;h����� G�l�d�`]EF�hw�զ�����w��̅�@v���"G.:sYBj������g��c��wo�"Nϟ<�5{ii�_T����p]a�HQMz�X��[�#��}w�m����V��>��+�o��#�:U>4{��?^��H<�]����G7����D4�#���&B�cڭU�T՞T^���/{��!��L'��]&͒G��}cB�Xg�m���os���+���6X���j��A_v98�\�yԶ�﫱ƻ'�bS�*W����0��O.�(��`5EО Ȧ��y��vh���BW~+U�E�E� �X�&��m&�#p��deb������D�"::��wgI��2MEf��o��^�ꐈƷ��,4�LM��b���iCU׾�:�$�2����#�H���hR\^N�YM��(���2�򁐑�]�oui�;N���z j��6D��\�дK[TY���>�u�09!%��_1.D}Ե��D���8��Jm�pݴ� �.��h���q����!P2<�;ʳ��m��L�,c�>R��3�T���y��z�I�&|�c[E��'s����$���I^η����e���n���{s6�}�c�.�LW�b�_�hkL��\������w�&��+8�IM/�U��Y��'��!K�C\SXG�ܒ�LJe|���	�S[�3� ��)����;�Ē<]7qnfY]z�UB}�LԼ\�<F� <�?���#��\�U�N��P�3C;X����%�E����� ���x�lhO����z�$\X>�_*��H���􉑺��9f&_߱@�^Z�e˒*�<���5�&�7~k�@��w�^s)�_�n}��dwh�����
�(&R���h5�����ZC���t�Tz��E�x_��C�j�J]\�d��i�Iٵ��˽� ]�����<P���pD��5V��~ń*�k'�{}����T���C^��yP8����j��Z\i�ޣ6+zltb��<�_��j����!�@�X���:�-_� �B���$�r�L��7�⫓�9Aϴ������Q��l�� ���H�Q�Qc��f���-U��(]�3K�������wn[�hʮ�T����O�䢫!rG��?�y�6����Ⴓ�z��Z�ImN�m�"���)bkN�=ө�ގ��%߃ۙ����k�s+����Kw��_trIn���L�fV���t��~���b��t�lI�,��9_b������ E���t:���_�mu+��p�vo(�cS��%*�D�Ţ����os��`w�}*{m���εo�������ػ�����CF���Χ�Y*�ݾ��͚Uf�h��>c_.Q���H>3�@�FB�y�7�a��^�
'FI+��̚y,EZ�>a�4�!5Eyd�5^X�+R�u����R�S�ٺ�n�.��ĸ��.��S��n@b���c(�ݝ�����k\=��|���m��M1.�����o�[�<�˜4st�nS�N�DWq��?���&wg;)W���
9�G�$o�2�)�[�s�z������_�����;y@��0�ߐ�W'��g�;?O�-߆��D�m�m�X�]�s�B��U��\�/G0�,�&���,�G�.ؾ�L?�N_��nלs7X�4d��h�Jp������v�7?>�ґ@4�����&��g��n��7X֟�}��X-��F�><�V�\�:��4D�/xD�?��2�vIg����X哴����������G�z@����Om�l�YM#6���)�%<��e�7���m��i�L�n��\2�;l�
���#����h�� ��E��*��3�X��3e
�<|�q*ѥ������"��F�D#��4�h�p��O0O�Ln��mVf���R��[J��e��U	=}Q|����?z�i9������/�<l�8�����`�o� j��OK=
�C~��gÞgC��$�2U��l�8H�/�����ܮ9+=\��~�V�zMv���4�����D�v)�]���j���Nx����)��[�3^�P,��`�X����
���Π���"E�I�Wq�Ƣmf���$	i���AW�]y�#&��<3�.;�'8`RgTE=����3U�"ijx<n���M�E�l�7�\2��&�dƒ�qV򓟞�u�d��n�Ada?,�����~s_S��Foӭ��V���D2}����p�:�W���%�[�I��B��Y
j��E.G�GγVF���慭�`���u��Q�M,2��C�Da�l�e+F�L�ax-m��B��D�cd��m��f�yS0���`�������3�c���F:���J��/��a!J��{';�T�g�ͧE�ǅԛ5��h�0������D�WM���/1���H;%�99F��#�1��i�E֩P҉sͪ��=G���y�����W��W����A�sQ2�����QO�vS�Qn�Ď��X�H����'F`Uf�����PuX����L3�T[*�m:�����+ȣ9ȳ��ƾ�˻������l�\�����#�d=W����.�5_���M�#u��9�����"hGr��C.���s������ZTN�>�x� �l]Qs�m�mv����؁�NU" �DN�x'�Q�#��>c7/`��%ϲ| s���^o�e���.͞b���n�~�ӧ��8�4�����<e����|^��1�qe�?�}x�qi!$�ř��Fa^��6,�p�Y�K9"w��Hĕh��h�l@��Ӏ�����&�Ͼ;�䙗n=�q�����ſN-��>� f���g�xv�>>옷�4�>u-:>����:�o7�Pj|��Zr�(�:Ak�F��Ks�[�ц��0kk�����^�&���V^�¿ƖG̫�Jw�Š�y~� 5����N�\wZT�g4\�[���!��#�\n���;AFF�賧��w�,��[��@74�뚷�>��IKۭ���tO[lI��Tǝ���:q��i��)�B��y�L��-F�.���>1Q����Ԉ�3#q���(�\��ȷ��k��:�t��+�l2H1�r��R��^�
=R���p.�>*�P��'4M�'3b�
�b��O�����{�+�	����w�f����� ��(�ն�f���Wh�9:�s!R���o����(P(���"�C��˸
��ܢ��Ew[�v�ao��Y�e�ϣ��G'�]�tvÑ�#?�[�1n1�]DEvr���c�:q����ӞRX�1��u��sy���͵1��7�	��!K?�\_��s�_s)�C��HK��x�am�{-sYZF|���K�Q��P�ӌ�����e����w`�Ӊ�_oF����@�և�"��8��^�-ϭ���5�(�t��Ɵ���J��ZT��a�ic�xaM�0�����r������h����	b�O�ubIb�S���.C�b�Ȅ}����?��!"e��� �
�W��,J'v��ȷd��Q�P�ڎސ�🪳��.V�Q�>,�BBh�'F��6��vձ������	�J��rB�Sgjk��G�����sE,}c��KKЃ��w�$�,�ϕ�/טBcJ��ٰ8Z��4V����n �ko��|l:Xp<غ�A�O摲��/�˕M8�e���s�6������<��b���^�����~"S�t�Y�;[:m�"�k�&���&����i����7E����,u�jci��R^�@��1ԗ��݇'���h��Pģ�{�M�+(($��$*(�S�k�n�ؓe�ř��"C0�X�<�D�S��������l�z`HV�+xZ�����x�LA)�j%���휖ǖ�٥�4��.z�Ƨ(/T�R�j��򈜄E�Y���c�YT8��:����''g3��Ȫ��a�����A��������~TM1���-�E�{���^T��R���"ɻ��2�5���v� D+���X
dlt��~I��\���G��lX�O��
���� thT�]��q�L�b�c��C�fF������{amEIf#��tY���>�|A����YT}(���7_@��H߬�)T�(^Ԙyi�	��ql��n�T����Z�8A��Q�f�&�%DEe�h�B��\��j ��ѳ��%�=�Avq||?��W�#1!��D+S��wĠ1e>�ķX��˹�>F�H���2K��W`��> �Vy���i��~��Dk��yM~�� :nx/ٹ}�IZ[����>�p�C<��Y/������2����j��K�ć����zR����-f:���+��F�,?�%"�F��Đ�!D�r�E���X��r�j���'�����Z�-�Z���	�͟X�E��8���.P{  b��Lc�/���NL��U&�����}ӊSN�e�䶚�\T� {U��H�v�A3=��\�4�JgΨB�9$�����/4��*M��#
m�a�{<���,�Xt�s�??#��2��0e�;�����A�� ���v䢳iw~ <���PT���Q������j��J���.�6sFc�i�_��W
�x���y��p�d	�C# e�7O3_�D�
jx���OmmU�%z�CE�LEu��Y���z���Z�����5����(�������=�m������'h�B_�a���*���f�b��ʔ�4�c��R�j���	D�o	��KV�о�Up��m/"Gpu�R����>�8Y��l�����e�"@��9dg�m��j ��\����9@��i��N�Kq��8w�IQA1~����q���������V22��dh�HC���G�1=��!Q�q�͟���KTS������#'Q㇋���"^�mI�>�+��6I���t����g�Ic�es
jC*��`���n��K����u�u��o���YB���2V���� �<%g��g�����ky���ͥ.FUl�U࿿e�с�a�`�&*9�q�2pB�cBd68 �X��B�UX;�S�u_�53��"W �鬍�4�f�����Nc����(3��[şO��0��BJ5�]\�a��X��R���ʸ�m��֢��A�ե��m���g��)v^A�ju
Bdt�o��8��k�N�[�.nnR;D<��̣WD@�$S��F�>P�K��ɦqb�
�f�?��iE���
-�\|�Q��e�XF�i�����'��ьY�Ɓ^�Q�8��.��P���*�5�N����W���WA��l��B���|�q�.:B��Γp��+�M�#�l���C�?U�;��W�3I�	���4�?����zL���Ա�}!���Hy��Ji����"�Yl���C��s/N�'��)kJO�-�#�a@�,Z��L%OĐqM�?9%ZīZ�H\�(v�Q| $,�@����R.�`��PRC���.�����=ZM�\1t6�� Ǵ� �amь#��X'�{8+n落Pm�[����	��	���j]GBF��+��4�p!4�U�_��̊�zw���8�r�c%61}+ɏ�+�c�*(𸂓�`�����K��R�H6
�XȮu�;L�@4&�2N��rM���7�>�gJ4��BKf��Q��<�On׳v�^�ߜ��)ѯ�
h�0�3;?:(����#��jm�+�9�dU!����ه�-̪b��6՞~���cn���e��E�lq��2��ZR�Ѝ[0Q�^"�m:gR���lE
��{�RI�����G��&���%��X4W�P�.�S��~�ѪK|�>��8�#gPgJ��<y�j���� 
�+�33��v�!ZLA!~�b�kvp�]���pL�.���e�$J�����ȵ �r�����Eq�;6v;��t��Y����,%�l� �u��Қ����V��FMb��r�t���'J;)D�1:]��_����:�m*ɳD<�����et(�~��*%�Ki�F{5�b�(�"�Ea$_���*�o1�͔TN|���
=�h���D�p�3�l��4/�a5�/�|��,��rz7v�4UOú�jv�ȥМ���0�zn�,l�t���!T2=P*G��9��~?��0�.T藬��j��7�gSL}l�D6���N�`Q�映�y�N����3~1쟜Y��6�o�^����3,w�}��عP�-w$J1��'�>�3�������������Z~GA���(� �w��22��c��d-��OZ2�������2�qHe8�%>�n4�^�l���MN�����F��Gp���''%3��Ζk�(��b����ȣ
��"D4ڴc�E?���Cb�ndR��fYCK��a"�q��%p:�0!F�a$F�e���h3\ݙ�Ç5��E�S>mt�O�K>Ve�����ݞ���n��1�!<�R��'unL^-��'I TN��ߧ+�ì���ZA�4^��q׍��󔚰.�*?���,�i�/ 3���Ts��2����5)1�\�vҒ�md�"(*�;D_�q@j&>��)��så���<<#��R[	��V�%�v Ќ鱷����u����2��1��2,4�V�`����b�n���`�I������ʴp��y<Dl	I	���.9�8I��W1��������W�m����>PP��f[j!�_�=/ȳ��ڲt^�\E�iK�P+n�߿5�u^�|�s)��&�8���L�D4~�Z�� ��4��As�L߮Rt|;���ɴ�n�h�=�)�/���(Z��3�o^S ޽
٪�V��[l;.���ۿt�	���ŧu���2�ۙ�hŰ������_��|s�
����g9!�X�_%�;��Ik}�S_����ޭ���O�b���{r��p��h�(�QN��D����>r�V3�6��#�Dc>5.�m������Of&�9ޖ�R�gk]a�a��Y�����hr�xxDq���űlV4=�w����%���u1n���kǧ�;&$]������B���r�c%����߾Y���|7t�}r?�_��%D^�
�}�
 =��>���A�Q��V�s��/��/����4�u��ԩe��I6VE�m=�:{֣��Xq^]n&��K�h�rR�{=�65�T�>����UX��L��$�g�
��S�� w��e�bmaг�vAB��}Y��-4�;�,_i8^~��D�����e��a��v�L[�jK�,�4_�y�GB�����3;�㜨�2U��l�t���/
��":������l��4Ȃ<5�:_�>���x�v���Z)�L��;O�|@m��Z�yѡ��qa�]�Ly�س����]�����y�I!���r������Q����;�6[����_i�0]r1�9};��e�ݻ'۱m<&�6%���ٟ'�@����Ş�T��SO�5�?�����t{�p�<S�v_4�Ob�u�e�p��s�浺��}�1N���w�/�xru? ���;��w���.�}�&�>���w���"�;{���r�K�����G��[��;u�����f�J��KDo��[_��f�*ӞF�qJ@e���U�ٵ�{��\�ϥ���L*�ț�5�	�!ε�2/���ӭ�Q/��F<�c�6"9������1"��"�PF�4v�4F#����9��.����z�Ͳ���kx���2EV�5�5v�fY��9]��X���������Z�D���������v�d�#��n�����g)K��~�_�����¤H�4pmԥh�g�X�+0��5��AH��3�Z�7��i;��Y�$ J��JԜ������y�rI#�l}�o��R\����8&�t�t�m;������ ᔌ�Q�>��ҞNE�^�H""���(�w/<<��[t%��SSK��.XԙF���߀o�e�/o������i�����:%8_��8t�9���Mw>��4vb���Ӗ_ׁ��pQ~�k~>KՅE{�����Ph�I���ڗF��7Ѵ4�琯	߹��c���N�>b�j�~V}����,m��?Q1��(Ҭ�D���XH¬�l�f�P�7��/�p2��Ӡ�>�i|��9k�z>��{���G�
T+[�ݭ��D�׉|=�5���9�=���8���7�.���&�(	�.X�ת���G%G��a<N�f�<���7���=��l�X�=���R�&F�\�Ph[)W�{�O.%
�Q���n��"KV�ro��ַ���@���2c=oO��A�G��3�����r{^<���:�_?�Q�h�F�?= �lAe�?��l���G�aɫ�Ia- ���[��k�dS�j��nF�1���W�N��^�~��m���������5��8b䶽�?�Yk�����'�M�n��bMcĉpq�8����\S��A)�['�SƷ��}���Jjr�FEc�k��$�Z��޳�Ve��nQ}�҇[��w�:)�G��d���Q����[��i�'�_8
:P��՘;.��.6��ڛ����\26�Y�7�hG����@!�~�`a��}	��E���_�L�#�dg�!ù���29NeVS:��Ebݼ=u|�uT�f���`&f�w<hd�Z��4#�lw���H\����ڳ��Q�������cbڟ	�[�y�^���R���)��î̓�@[���ս��p3tg��'��\���'��V]_tA+�ռ��̚(�!�wK����7u�uL;͗�g�0�{e�� /����J ���(D���i����(�Č+ׂ�'|����H�ᮄ����p�(?#���׶��:����f/*�� ��>z�|�|���y�9",mW-��]��b|u:���F����^u��`��;H�`zPQ�[�:"�K*K>;�!;��_���-��6&�g�[ʐ011�ǰ�G yj�a*|)M��ڀ,��,��Ǹ�0LE�t�X���EҊo<�6$v�<�zQ8�i�l��9�%�w��Z���fuJ)|j�&NYr��*u��%@G5��0r'w�8?ry]�z��h ��B���h�d�pD�j4��g��`�;���\��0o�Y)
5�l���<CeW�����8͊l�"�z�?&��(�>�5�C�F�V<X.?���Y����ew\v�p]z�~�3�����P����:`iե0w*��Vyں֐�~ȍvz��]���qo5Ż n?�������u��!�����=O	�/�{�Y�;ޫ4h
-6�7yd���$���f�N�D�����G��u P���W��\����Ի�}q&^
ڌ����?�S����G��SW�0�� ��YC�\�i��^��qO36�C��Z�qCkPL󔛃!>O�jf ���|`c��Z8��e{" r8����F-a:�u�8�oΆ@���+#L�~�d�ҩ��V�@�2 Z\i��ЛC�ˢsY�JSc�x�oN���!�@��K�L.��ʒE6�'�΢�ƺj����ݬ�C��˫�F�t{����<E�&�}ا)��K-#_�X��Ìff|܇V�l�\d3��!�\��#_b����,%�̈́�+EZ�5�rx�Ӑjt=a�(����7�������4e�r�*�(
]���R�иZnPD:�)����e\8>��07뒱�A�ϔr�"���\��hk��~^h ���<�Hw<���>^-��)9c������L�����'�e�;�J�k�T�e��	���p�n�d��x�y;py`6&���1XD�NР��ҵ���]������
׹Q�c�u�|�rJL��������1K.�yH�S,�-������z���7{������H11�8��a�]������q��r�t@J1���m��β�t_Lb�B��*O&��G���Vh t��6'L7�K�<#Qr�����:����%'ǅ&f=X�9�髾G���\!+�Cy�pm�ks�� �<˴�А|-X�cvq>A^ii­=�t)Y��������sW66���8S�5:f��#��C��Q�v,�!Iӥ���q��\j�J�]�s"��Q��t�J�:7e��$���w����I��qS���sMxF�Np�{DCl`�-^+�j8�c�p���7S/]�y8�3����S���8)�(�o�.F�(�Xse���A���>5g�$����:��T�������n�G�Y�W)�d�΢�`���b֟�����J)����BN;��l�A�9�F��/��)��앁�y���S�����;������׏��j3��ĵ\2�9�(���@�=���t���u]�xb�����m۞ض���ļ�Ķm3o������k�^�{u��v��ǸG��YoEj-�,�O���m?�L�m����>(1�H�.���-2pɒ�tx����[8�I�k�H�PH8ٿl��fs���Map����+P�G���uFiw���`�ɵ�)}&D��M�[����zO�Äz>W6>!Aʯ�e���l�>v���r�Q�X	�H�J-�,�ˁҿ��6��3Tcک��X W�L�H�"���,V���}�	~��}�;�A������.gL_�$L�kK/���g��8'�9���*���cI'�7������.2#��z �o�N�t�y-$��b^��%��k�s�����	>t�=��S3P�+��r��U��Dl�\�d�O4<�޽% ����q����?�Z�]����&Ъk-�G0�q��C/��H��d������W�c��;����t��e�����v��
K�\4h:�℄0���H/��%v��e�V�������po8�B�����S�5�����T��V>)�4�چ��K$�2�R�[k�^�֦�HE�nq����M0�8?�d��9�A}L�R*�=-��֫���q�~U߯e>���_���٪{�_bX�kc��HD�[�;GE�xC�����%��ZMN�iPi�x�}�j�����k7����n\\r.�ԖlJ���5R����e�? 
�!��Բ��p�+ҸٍЪ+�J�)����۹Gl�Id����.IH�{��C�����1Li�L�xfV�H�� XA/��*ZAa�&����ёp�E��}�!o��f~s�o�.�v��'���"u\T�;�7$h$���Ԓ��$�i�4��7�4�|��von��+��&�D"S(�RU�Q���/Y��?��"Ъ	8`��O��N9�-W���ܮ��a���Z��N�1����"\Pf0�����P�,����tU�U�U��2��4#�W>ym��G�GS;L���/�Veͽs����N5J�A�l=|F��[h����l�Z/�N`�)�d=I�Dc���=�Z�5[���K֚��^�ǖ��<�[Qr��3tb�I���pM�b�n�*N5A�ISS� �I��"ؠ)�hD>^���\M�9��X�_K��z�Z��3(;�9��AX$�1ܭE���3�s�Y"��{1=`O��]���'Q�C�ґ�"���bT5u��_��H<a/8�d�o]=�� O��{�����O���1riӍ.M��o�2J\ .Cxݗ�r����tz�r��|�Edm,�vC�ē�
c�w_��z�H�^�,�\ȷ�N�+�hhڼ؜v�pzZ�r�EUb��*�E�*���	?��9�-��t�V�)W.��D�o ��r�mp�@$7���w=�
xD1���/X�\�+g#Gn�I@���ĭ��.����_��㜯i?�'[{7:�N��Tq����Ӽ��[���H �Av����g)��-a��,��V��)8��|��y}f����ԁ�2�LT%��A ���3���	��E�}9��e1�4�$�d& ,�&��T6I����>�Z�ȍah����z[W��r���ףʭ!��D�P`|BpiN�,���σ��n��'-K�82�-���	v��0'E��:�@*���F!{I�5�t{��Ԅb����ְ&���[��d]��ɘ������}e?�v���F��ځ<uM��D�:F��VU*��E‬��������0(�B7L<,���.��3�`����`��k�D�Y�C�]zx���G<(	H�,����`R���tm?�5h�*�SGe���kQ8,�t�� �\Rd�.�b�A���,L(R�^lH}�M�~[��e)t��'?�T�n�Ь�]�&r��њ�6�WTD �}���N�*g���Ά�b<�Y�h��`xxR5� ����%yw�ErnS��Տ�h��IWF}N��i&�V�!1f�̘n��M�X�IpM:��������`�pbM�d50ɤ1����&�{��//^4��ǻ����<��id�=�Ny0F[���D+�;:L�Ce"i�[�)����2�+)��$J�(� W[4�������:2݅� ����7@��LdIϰ<�����Y��7�h��LY�Q�&��Ux]v=�x/[Ċ�_���*��	Wn���u�9��9�i"���Y�Jʪ6��G�dk�+Ѱ���`\X�2,7��<@��YI�0Z9Ms��!?)�VC�WKWD�n�B\�G��3?Z�mc2l�jc���K���KʝH�2M�����L [[�.��]MG�1��f_��lR4%����~/�����IIQ5�I�y��js{��ʁu�5��6$ZWQ�����2�00n��x�ų�󝓭aw�@��lo�ο
��L����*�Ag�1nQ�?�#��� �d�#��֏�g�y��X�g��F����ㄔ�����L�H��R-iEZ\��� {ү�"�_��܆y�Y���
1vI�r��!@0�(ϙd&#;W��E@��M�Bs�R�]e�f����m��-���O,y�'	�\�G�M��d�<�Vsj*؊��֖�K�������~���a-Wä����3+I��G�����_�MF�O�{��[p'凡��	4hiM�}�q��Y��9�=����t�a�R{G���N
�y���r�65Z��L]�N&��g����	^u<��\�DM�~�[�z��F���q���~�W�nv[C3���R��I`K�ggc�9Z�D�m>��[��s�g\{�8k�9!*}{���l�b`0���+1I%⻏����X�k�ɺ�H	�J�����ERF��?={9�*k&N�yd*����_	��U�����Ԕ4��I��x`�g�Y���`WeY&�Eܡ:=�鎜-*�ޗi��A��3��ZTD9�xP�t>�ʝ��0>��٣C���{���G�px���E���)�bDA��. �n���-�wWt3�%@���oW��Q]x��	;�u��)����1��Va���]��7;��D�� "Ǎ?+�=-���2i����K��^ۗ��OxY�7gD��e
#G�P�^���_ۡc��,���;C�2���
9����2G������٧qڙ� ���������'�Sk듫K��ɹ�9�Q��
��T��!0,����!Ek�}_��z�/���J��ϠNMg�+��p��+���p���ey[�d��+�[`Bu���,Ap�a�7c�˾��M��ݖg2\�+{'&cʄZJ��0�f�U�G4@���tm��aL�{ހ�s1�1��̊�s�]{�zk�
H#ff�D�N�b���h��%�)�Bf
���0��tzϠ���>�E�A��2d�����%��쁾d^��J���,vpw&��$�8��ѓFx��yG�`�0��Q�<ʚr�R���""�����U���%�Pm��K��ܪ��p��}޼�6����/�Q3z�rgO��f��(��u�6�֮�,��p [�1uH�>�L�f�#��)��
Y�}�(�Ɉ 8����Lu����r���գ=��(�k��װx�y#G�2�%>�g⍺�ĊMD3�������U �D��Tf�F�7�q��������)6w���3�U��{������O#����"����m��W�e#ż�Gs�m������|�����,&�=ڕ���ཞ�KT^߲T�V�ۢ��_��(���,��l�!�~UI?��m�7^v�M�,M��nI�|����ڰAq|,;ˉX�p���w���'MF�}�et�H�0|f`��C����\�1@�
Y!߬;�߄&he7ߢ�'g��n/��j@���7.qK�M��;6�A����o���K������֑<~QOu��ם{��#�[}��$?���X^ˏ�,$���_���ui��!�/8S�v����q� X�X|#oJ�n�?�%�)���>b��SfM�l~����%���6�PM0��� �1?��zC�ؒ.HN��E[Ogj�}<�n.��.w��Q�k�[=�6s�ߴ�~kx�]&���H`�+ug
��	��#A�!j̎��,o� R ���o������kr~�p@��
X�R����T]?ŖSWg�l7���w��}m�#� x���=��/�_
(���S�����{"������4��1Ĭ�[�F����y�L�P"�\2�7b��G�Ǥ�K�)�YH��4�T7'\M1��<�0
����y������6h�����?�l5E�F$�g�{���ܔ��!N	�J�x&"zFn^��a��q�L@;���4^�����`���hݒr��A�֖(4�e�J���Q{iv��X*q��pآ&�j9��#�����|vZ��*U^�R��.�H QvSI�Nȉ�TSXP��>���^��s��m
����h��#��D�2���I�x�"A�'ƎCU��=G����_��F�ٿ8W�X(�
�(T'�)�e��HA�])]jfU�?{O�>5���H;�J%��P��/9��bE�οs<����U8_�˟vb�#�G��N��C�^'{���)�n�
&^E"�oW��7��w�D�Q��M�`�6�"R�j�d�o�NCcF����ԩ��)�����4���{繭���Ʋ��xl�{DN'PH8�`���a��<���/vC|ᡠL 3כ��ڴpO���HB�'��ң���l9�����ħ�)tpu1�rs\b����N�O2Sa���3S��y���Z���?F��"e�c��8gu弍�ɣ�fW及�w�9�OE"�Na�]�K��[�e�^�츰�w�Z�m���l�$Z�T�w$9R��8��`���9�~��ၖ�9�$BO��\�F��s4��Ƥ,驧��\7$kW|.kr֌�� U{,p��ބO��$�=���L�>\c� �r|�Wq	����uX�I�~�ƉT����.G�,))o	z�� ���[�³ɮ'aPL�C!<22�I�����~i�%E��F%Ͳ�	��~ˠ�>ݹ�ɐ�B�sǊA�'�1_��l��z4��VYa�Ѳ���uĈ�Tl�~��bS�82̳C��FkXD��������X�����Y����2�^��0j�Vo�p�P8�F�9��5=�S�hg$9"�gf�Q��n[�ߛ[�9��Zc�vx1G��X�B��:�^�,<}�TI����V�bv��]=�b�G��Ka��I>�X�G���?����;��jl1��i��gRx�༖+Ҝq�}7�^ߑ��K �֋6�?�Y�|�~�l��t���_�̘0�Kb�L���+��x�dʖ�j�8%a�T4�葞N���r��BC6�a�:��}�u�p豧KM{��t�3
ǭF̝������^�p�LC���qp��f��Gb�j~��S�Lg�`��H-��c���D��Ə]�{���1�p�c p�ޠ1��R>��`�l��#�\���ص�������c�6��c�TUU�}NP��(�e�F7�C.l��FӇ��`ڈ�F�#;���ڞX�'��a"���*oS�Ǻ4��_�6�T�zJ�e�T�p��I�+l���;�_;�Os����C>B�����wF�&(�0g��2f�z�FI/[�:��u�]`����H�P}Q�^�H����;,@Ow/X����T.�R���@���1�E�qx���|Y���H����Sj/Ez�,����_	P
v�)NA�/Œ�"1�NZ4�KhVt�D1l%ZO9\m)���۫J�����b�P�����0dTD��  0v,|pM|g�۽�t�<�l)��$�&�ܛ?fW6#����W״�5@�k�q-�f���n%�5���f�v22ڬն :��_�U���Iu����J���d���Է�Z�MY[1�jP6�o�	���J�@Y2c�h�Vo��d&N� |��G��@+y��ڄAk��Y�Q�G܂MJK�n\87:	���/X�.i:�XV�����4���*�y������ħ�̟�� ]�k�Y\���Ʉ�^�/g������M�8��Z_� ���4��2�B��LPM���0☀U ����*���n��Q]�M�7�H�6Wt5�-.��<]�ČRS^H��?�J)i6|��4�#=j�"��.�X�������6>sS ��z�ߐ����ꀆ
�Q[4��:����8�|�����`h�_��6nJ/�r�SM�8��v����Q�@N��SE��1�u�t~����'D�ϲ��Jc �F�����Q1MN-U�ww��_�Q��K�Sւ�]bڗ~ֱ���)�͐ۇ��2�W[��Dg^�ԩwi�"�-�J�	�1�(�O�U7b� �5" � ���n��Ԛ��4A"T�l��G���/��z���^����~kVS�p�8���&	���&���]t�iW��b&�QVɚ/���c}�:����&VY��6>y��s�"�8Y氵3��='�t&C	$"�<<c�%��_ܬ,�-�oEC�����8xE$Z1�'��5Ml	���gge4:a�J'ܾ�?��kk"�����f�ޥ�G���S����NI�
T�:�9S�py�4;��x�U���W��c�,r�bۧ�E�>�R���zz�C6x�w[ێ-,��Kd\����n�����M���0ܒbl8$�~hM�͝�R+�u��#̨R&џj�3xy�ݼY��B�ЍcdI&1�@�*��:��Ĕ��j��ֶԸ$��������5�5y���ޗ3��R�z����X\%�'5F��4	��Nt�о�6Bh�'[����#����5��$���-u!#6!�ڱ��|4ݢt9CT��@
�&�*�ESM@A�P�����O�irq�P�KC��<#W�DK(��6>�G�-1gcR�H��vY6�(��N�l����J��
yD+	���*�.��oU�|���f}(]X��a�&-bL�G)���yW�0]�?���o2�����u�F��N��{ם�����ݯ�es�ª������Gӡ/xW(�b;j^�h�c����i��lo�>F��%��]��7�R�n�]�K�է�	�%���1W�<�9�X�.�;@�����yQ�%����t׷�Q��>���(i�ִ�rQ�[�-K�z|��~#H��XI�(j�@�Q�%�\�W��f�M�)���1',�*�W������g��ۥp�D��.q\��o�l7�d�e�>oR8�����Gp ݟ��5'�PHik����[��%H��S�Gl#/7�����ŉ���0�q
b��QH%X;��Nr��R�-��2��l��ʶd�ڮH�����ʙ�D����lW�}���skkkk6�!�'P͛M���b�W����v��Q �7�g�RN;\�s˺�ʧ�e��U�2F��X�$ȿg�8AȨԸ ��!7B��3�7jR�ؤ������nsfT�aכ�q��ԓ5�6 �-��s⻴���#A�	�e�����wE������%�?N����G�S�y�]�VeuFr��wD����t9�eP�i��n	��q<ҽ�d	w�;�sO�u�
�qdh��o+�ړ�G��kOI���5i�n���
�ߘ�h�%��}�������&a܆|�XSN�Ǣ�'��@ 	@-d����L/J�`�b����7w�����_*�g-]��2x���r�K�KȤZ�1g���=-�x������j5&��[C�����3�e�U����v~x����P��3;�lqֆ�)]G"W�ih�a�D=�9{��a�e\9�)���33�ڒ�D�og�U����J�JY���f�����4�mC�l�	�����?X9�J{܉���)�G)��!�k�ٻ��4b��S=� ���������X��_� �]�����P�pyI���{��I�8�,���ϣ*����l>�P8sy�6�
:�(s����e����9N|Jk�y&;���`����_�"�d��U���hfs�+�3��"�Z����L�<k��OhDǤ���b�Gnh�#�W�l;�'����y��1?��n�"ǆW������*��L��G���f�-�Pܶ��J�92r�	��������E�����~S�M�B6�a~����s!7�WO����k�Z=��4���������u�����>���+�����E0��}/�����yі�b�e��~�~fjUˬ��	�u'&���h��_.h%�7���>�/�Z-*���0���]�=��#��z�3Ѻħ�����n��\"3�{:��z�P�<���R�ؠtS)���v)RZ�'����+���N�D�jD����aݡӹAͶ���o�H}`�k�,���=�f|5�כ?��|U�3���ep�fqΟ��>?l�ª�U�����
�2�ґ�!IX�h������3�	�zE���޼�CLZ��VS��H&�=�z;��	k��[-+�DΞ!\��Q8F:r A���">w'���%��;Δ���㛽�T���3��������vJK������ *�0ׇ�c����牡|W�#�Dhʙ���[�[���~E�����H����]�����惟[6������|��I *�X��!}��4f�
VА?}�Ha�a*��V�&e��!����"��e踕KAy�G�B����*A�9�Nl>1@�E(J�|֘1�b:k��DՍ�^7sγ��Rz{�g�~�8��m��9|�>`R>)m�:��g��1s�?�|�����c��z�M�����0�Kob���7v�K�s�_���KQ}�*��vo�^6�t��c���X||�Y�4 ����;2W-���/�j�D�+l-򁅑��i�~h#w��lC��7���ں���J�x���tZm��lZ�x����w�dm�	���̅�מ���?u��y��
6ޤ��e{��"#{<��2������D|���x��(�߶��<���-���E��g����P�*��-�q�<�(���FQU6��.����ksD���;ܰ�ڑ��4��Eκ��mY�|���>��^i����.��[�/S_��g�w=��?}F؏��8�2	,@��2�U��#'��Ӻ�.�l��K��nG~۾2�o�r򔩲Px��Ij]�9:_c
7;aM%)˃�N�	��С	�jY1��j�,a8osj�&g�߷����n�z�pfa���Q#���t����#-��5H�Ԫ����g�Z.��t���7��b�ds|��y�b[O�n����Kvu۝�\t�����2_�NWy5�0(6���(�	�D���js`���>o&�p��lt��~]�p�z%P���6�ۥ;�j�R��O��{$6�����S&��>����u?!�l��V�0����8}�� p��Ah_}/=�P�:ш�3Z*"5�H�
�Kf�u"�IflI��ua]�S�w'
�m�	���g�d$�*�+�8ϗH�X��� �<��}��
�̚$#��IE��d����8]����ȽD��~SJ��k�^�r��!a)(�eڳ ������� �e�	�$���(q����\Ѱ/��vs���ｹv����qޟ����y�3��D���lџ�z(>|.�l.Y��ʥ��������ь��C̖�5I11Ȥ�̡u��yŭ�Ϗ�j��	t�*�j�������bwG*hQcD0���A
��O�h7�5��2F�Rͷ��2���AH]Q�q>�6����4��z�+����5��Rr5��?���i<p��y�RP>�/t$<�|���o��q�,�zq�k�WH퀡6jgGH>�/BwҳD%�R�zeG��Z� x�"u�ދ�#�!�IB�����wg�F������L�ǉ|Xԝ섉�q>��J0��0��Ò��KJ�h>J��=퐾����H��"���`5���#,Ճi����dՔ+3p1��r��k�JM����.�Ki�>��!�7���W%�+zP�4r���S"V9�L�����_r�6��:�KP��=5ɬ��7�0������=	1�KJ�*2M-�r���h�z���VS�cwpX�h���ty� T{_k4��w��f��L�$�;,E��6j�:+�G(]kn����H��S2T׼��s�=p��_�k�	*\�m<��c�2{���{S��Z0��$��ua��D����⹺ay	D�H��0H�h�0e3~���ȉ��]�F���*y�׻�E�ͦ9J����%���-aˑủ]�{�8�I��T'>1}}�����]ǯ�l���5*M��1{@��sVA�=m��mX���g__�?���)I+]��6�q��EQ2�a�0	'ʸq�N��V$5���om�X�n����Z7�{��ʲ�}^���]d����^�׺����J����.ϚXkO�{	���
�"*f^�=܌gҌW]k~��7�ц�S�J�R��9��E-2��a�r%b�����oPc�J��_�"�OM�\+ˣ�g�]��Ӫ��H�7]ii�&Gt%���r�|�c���l��0�|�5�2�ҝ�����wR�2"d�KQ�pZTk�arF�r3���?��Jˁ�.�b;�n�ʈ��	�VBX��!]�/4��s)�;�jsC\	�V�׭�|/�	?�cS��q8���BҮ�[��!�㯏��Ms�%c.��x%!�ӹd}�*'�h�m�0�lBqT�L<m�0���{�`0�{#¬Bc���e)	�r�]����>"�(z��p+|���`Ɂ������:;���`:�&gvTd/��rnO7uu�iN��r�1�Y����{�����jS���A]]V%MA�bA�������=9湞�����m�%�|l�)�o�2�v6F��]u̳�Z��q�#=� ��L�,Uڥ"�謅�Ň��9Y��;p�9H��_l�8�����ǐ�9<��2���I�4Q�����;�L]�j�Rz�y*�?C.�/���~V��a_������/Ty!�ѶA�k������[�������D'�s�آ8NICz�.�o�#�0Q��A<�l�٭�ǽ�{ާBgȒiB���6�&���ô��w$n�`{7���Y��H0Md)%����u��O�Y�&�	ʶ$N诨L�xu��[�����nxǲVt�Un1���YSn;6~-t�І�{>�
"��ݦ�Ǫ��Y��˔Y٘�>K��6�iQ��.�𽼍� ��V�5�W�'��[����� �˞dN�b�*�+��J�v>^	���]亸� �����fG'ǒ�]�*t$H�D��
�w�1�&3r/Js���-��]E�h�Kk�cX-Տ��G@��(��fQ��:��Rt݁i��;���5�?�\�`-�,yˎ+�ȓJrYmi������{�v<�����_�ToR���(	��>+EM�dQ���DN]<:T�B-D/���]�f�&��~ZS��V��)�~���a.�2dhnQ�O�)�N�9�b��d��Uh��;:��B��m�d^�`�\���ƄF)O�0�pu�mU+���Q�)���z�Õ��'�|��n�@���]Πo.��'��-`�
3�����v�����*�Q����������_9lkc4�����7�H�w��q������L��Z���1k��	rX'ujQm*�����p�ԗv�n�HK�N���$� xĸ�׏biHL��R�,��{©>�C}6 j�.�CRO��i���S�[�^u2�T���*�]>��2��v�Ē*7Mnh��罴�<��0��!�eN�43��q��s|w���և�<aU;:+gZ|�l�.�-^M=�h���������!C����d�,�n���%oL�aˤ�V��SЈ����\A��A[�=#;S�V*��u)j�d{&������C�Ӱ@��X�񌂯���4�x} �ҘP�:�<R��q��^KRW7��l��`����Ѯ'�<�?�#��lˋ7��#�l8Ց�N�M1��������mnv��pv->�#x$�6�-�����M�c���v�2�/�����s�$CƑ��&��vqjT#���H�蜃�>G�YX�9�>���I���0c�;"K�l�U�3wj���.&�g��(~b<6HJ���y��SWI)
��y�J�n[�*��HE|�Y���}�����a�:��7��c8��0���Gɤ>Mq
���=L�3fH�A,�_{.)���O�U2TX,�Q+4�L{��+�-<�a�Bo�4���iy`�T �^�|�|��dr����j��0y�\%�@�l���nɭHP�ds��=�*������qRTd��2kS���6�h��%�t@��[c�_�A�D�\�,wX��=4����V��� �(���&,-�ˊ�c�+�T��,cX���~hO*�\�:v�'O*>JҎ���x񮱃�sW&��1�R��·���f��wkB&�%���5�:t��:��ZJGJ�юS�
�un�:�����R��i�ҦX����F�S(���[��O_�Q�>���3(>G���(���YSr�	?�
� �EI���ӵ���ܲ���`q�Q	�T��XX�X$ ��O�P��O�7hT�i�D��\0E�]P� ��F$͆�v�KkB	:[�*jKHPM����Y�_Cr��.�+�RF�D����f�dxNO��L2�7^�L��.��R��6��Ϯ7���X@k��i}��# ����u�ϕ�P���h1��R�^��-��'�	;p�qL�+ÌI4l7s󦃭�jl�]�kwY��|'��""�L8k����-�F��FVi�-5��GUH��#��C��I�*�/�st6%�KŐ���*�����aI���Rg���[%�p9�řx�=�;����=@��2j���ǅT��/� ����)r�MD%wi����>�d� ���(±8�*�k�X9�IC��
�X�/@G'�G���j��sA�Ż$�x���KkJX_�da�|�YF�:#[~�j�LU������'�-E��6�T:}��:�lfU�.UW��<���	�|eڑP5:�o���Z{s���TTA�Wmqi�O\nY1+���U������V�4�ni�;n=|t��E8ʊ�u�U(���g���D=~�p�n\Q�8Q����#�A�摾!�O���)ܽ'�0o��}Q�Kf#(;s)�޽¢%����!`��Ƞy�Ƨs�W		\
��I�jq>�;H�j��?R_[��,	6vϋ�Q���z��0���1ש�O�Xb�'�4�EB��rJc�NH?D�2�Y�Vm5���2)�6������` |Х5#����rC�%��X����f��X�##s�Q`èqc�,r�O�Y�=η/]vC�e��ܔ��Z�z��eJ�6e��P6z�(���Hu� ���ͮwK�k��r���087�������c�l��M;���-T�,��4�k\`O��+���>�.�ub���Af%9O�M|6[��Fqxf7)���8L��@��+�yB5��As;m����<��N�3�Ye~�:=>���)���)��,Րէ�(���Ώ-"����@�G�+T��, �
@t��9`��ذ��|L%�\�a�<��Yo���UW����O��]��Z|V����Wu3b%hg��eЃ�M���Ν
2��m���s6��uq�qph�&�Z�i>|z�EY��j��N8S�瞑{:���b!D�9}�xLxUT�pR�#\6+B�����Ӗ�R(p����{�`���d��^��tTAű������*�Kz��k���즸QG��˚��	�w�I�jK_�M�	���M]�
h<�_>�����I�7�k�{�����a��7q��5����D=���]C$X{"��Ko���"����J�%ޭ��O����-S��7��]8�ċRv�`U%ze�\�|*a�@�b]����h�"�U�Bv�HHF�����m�@��:�4
�H������V��{{����,O���1�=7Dn&�C��M����N��T�[ݼ<��o�xf\�E���nC[vUW�<Z�o�$(Y�Y5BzT���&�,8Bf� iq҇\dV|����T�6f�.I!�vf@H�i���"�0�x@wg��4�����Cù{o��9(P�e����()d��2_�b��Q�ʵ.�6�a��^?q6k43*\@�i�D<��b� �h�ڝ�gX4�䡿�^E��2��kf�\�?�(�xl#Nuy����5��eJ�&� 9�|x+��tH/Љ/*Z�^aTy�}3��o�<V���d���\8{���?��o����� �I�3a^�a�4�C������X*��<E���A����!m�����~DuoL(cC�)�6��\(#�@݃jDW��#q�e�ke��D�d�g,��᱕~U�� �����J�p�rF���h�\�F��`��f/G�*Ɏ����.2���p_ﶃz[6��� *o"���XN�^������*�9�����q�yϻ,�
3o�>��:Pd�d/yDڣ`3�ց��
�CV�]���v��uKm���
f����iږ9�9y�rt�������Q���o��2�cB��lH)���|�KN-��j��!?�N�h�ؑX�z��%���	�o�J>���?�T#��������teq���Ɵ-��fs���$6?���#�+ 2��=�ne�W�F���x��Ƙ�6	�@�B�cX��� 1����耆Ɩ/;��2A��]W�ι�B����+D��ؘ`I����]�m-_v6��J�����ķ�E�	N�?p�z�N��E�E"�~ݢ=���p�����f��U�J��1����.��=Y��G�������ZqXeL�j�:�X3Ʈ�/+H%
w��PAi���ތ�#qu�o�Ez�t4TF 
̃�+߸�	5G�m#�1����ʼ�m�ѧ�����z�ԙ�FKX5��(��C hhӽ\�Z��O+��>�_5������:T�l܄K��G��t2�Tn���_�g� �b��`�|Q�'��������Ǹ�0D�%�$����1�6��N�:`���r�	����-�IL�Z��9�o� ���~���
��{�/�T桶%�ib�S&1nIt�p��v��]_`)dΐ�R���Ŋ�U��;tf�[2f2�AgNc��ʬa�iL��y���{|hR���=x�I1X�o�n��_T�J�͡��CE�|�{�>�E� �<��KH��D�o�G�	D3'ѯ�5SA��[Bz[S"}^�m�ݮM����T {,�`;�i�o�Sg@a���ԕu1:���҉i�Ǜ��nGL����P���[��O��X��<����ݲ8����C�K���#�'Ƨ'����W�Ҙ�Q�4dX����[Ԉ`�5ˈ?J�im�[��r�;wmHH�[��'#�HLř�.�9���p�(��@?S���׶}���O%$I8�u.-H]H�KQ�L��-����}������#_?�տkU��CI��|�"��%5�) )S�f���}�d�@�Whh��>�z�����ɻ̙}� v�g�'w����0�3J�%U{� �O�D�b�sߚv��: �ö�j��{�Nhr*�*M$0�G�-��3}�|��s��4�
Y�Ԭ�A#��I�bc��p�5d�零�U�>�CIm��t�3����g�Q�솏��CLt��@��Ғt�9��&@����{@��ʱ����v�^��)��mu)}�O�0���+ɷ�(�i��ġg|�
 �q��n��'4
� �����\�]��y��^�޲wM�!��� B�X��8ڇ+��i�eő���;cgS7����-���L5��Ѥ�٥ESS��,�l�p�}o �ӟ����E�!�h	Y�vn ��
�&�[�G!��+��։�czJ�#��Qm�0�X*�iٹ+�K���i_R�^:���V���*��B�����"��:�
0u�lauy�c3g��VQF0a�Y��k����3{s(���\<`��s�Hq�����!��A�}!���_�1@�}�C�]�;o}a�m�܋驴�����k��M�=7�j竑J��+��&��E�v�Wl�ݹPu��(}����
z�*�[����L+ە��2|�m�al0?>B�1����o��(�Ud9��)s)�$@Mq�����13{`Ĥ���]PY��0b%��Q*p���#M�*�I"�Q�?�K���}o�Kԡ���'_��n�~�Ź(�\1�9k��H�H��l5��U��*tQr:�rM���ĿD��`XBBa�C�>{p8$�6 �c|���U��_�%�֓��	f�K�׊F{���7Z�l��w]���&i�ضm''�m�67��ضm�Ol����qǸ?�a��3��{�\�f�iY����L�&��OP�O(Ѫ���39�I�,Y��)� TCՊ�0n\n����|�G��<�{uJM�|��!}��'��f罌���?�t2�u�U��%�L�W7��V!�L�,�$�ǬO:��y�q��r��uPY�<6���e3}��F��$���w�'l��LD������R�Yq��]���Bܱ��
��	��=>���X�M��5* @��qX�9�5)��3��%E!">O�����_0�7�Y�_�O�P�޻9V�%�(�������M�k0�%'$M^nv^se��>+�%�,q�����Ǥ�A{��҄��D�V�])�%��ȏ�-R䘛�h������?Ut%��c��6�S���	����M;�إ�$�D����<�Т�k`�D�X�HJ�;�ֳ�$�XE��T˖_���6T-4���!?11�2Z�7|�Y)�k��=�&FSu�P]���*����!t�������U�!iaS��
lX��L�Tb~E�@ǫ̓��3o���Q�K8�������	�~@�ߑ�PIM`5�g�)��[�w�پy��9���r�"W,z�����\��ݚ��|˹jlh�v�Kkq����CVY���:d؊��cu�޳���˭W�n�ohP�q�٩f�+�)nk͞2�8n�݌^���O�SHD�����}foaR�۾�{V�K��?A*��6��D��٢r\.����	@�Ǯ��+��T��0jQ��i��%vP��L�hgmi�rZ����qG�FZF^�yn:I�60�?�"�bAH��Y�?���-$���
,`��>����_�U�._��QiRQ�d%
�r��${��e�٬첥���ORTA��Z(�6�&���`Äz�>#�ֹA}h.�H��u��ޕ�2�9�~�.�!y��g��V�>|D5;e~~<o�ٚ��K#��n�8���-Ϡ��$��{}}=�?�'QW�����tւM ��L��z1��g$[�@5~�)� ����=��pbCbX��'HZ�\t>)���ot�DGˎpĚm�ʙ�0�-��Wm�F����5j>���K=1[�z
p����)	�"]\Top�$�R���h䪡^�F���'���)��v�:��Xuo�À�E���d��m�䏌b��#�����b�FP���6��|���$jȊ����-u��'E�;�������K���1Q��J���<5q�-bǑ[I-Fs1q@]�I�ȩ$��@=b|��"��\�C�#)#ݚVT؈zw`������ew�k"JK�`��lEIMWx:����62R�ͧ���i�d�x�5�~Ӷs���� �AG�szz�9��E_�;����&LX����,���P��A|��$`վ����y�-�N�Ӵ��*h���m�+u6��l����ڬ�C��$�R%D信�Q�>Sȯ�B�U�%g\������u�޼"v����l2h�a5����&�����k&`AE�%Ct���ڲ����c~
Ȋ@?\����⬙Zi�ڧ�ן�QB{*S����?��}O��%�G���߈j�.Pw�=����k+���=>>�����8��$����M���+/D�(s�8��s�� F���.G����ȕ�R?]h�N~�OY���2�{��(X�5$�c�@��[����|���9Mb`ɩ&��nOHСUU �(AB�������e�ln�����������4e���+�촱)�^;d�qWx0�Ijv���#s�l��qGG"�h�`89%��T��w{3t������j���=�סl���P�צ7ϣ��{�R�sI-X~�@�4	o�e�c�wgѮ�#i@F1TB2�fz����\X��/�V������-�m�hP�����ON$��es���'��0�\os�j��B�.��Ǘ���=�����;τ�jl�EM����B𡙑�d���	�P�`���X��|C���i��i凤w�|��y�
"��8�$L-`�tb�����<����͟����\�yWR�l��16���z{�*�K� ��/���
9�����3b�4w����Y�{*wg����o�o
G�Teܵ�߶�~�7����w^u�x�3�Rp�8��6�ә���-�	-����Tc��p$��r(+&��)j5:�s�x��M�󺏟���Pp��	Z�0;/����W�]�WK�[��I���AВc��W�|r5z�$e8�7v�r�l����"��Gi=\�V���Q!]T����� }�K��>�ӂ�'�NQ �߾��k��E���G�����������b��m�HB�����-�*"ת��/�x\Bw�S�%I��xӖ���hK�"���6'�ʗ��k��C��A�)��!�(A���.�R�`�)�,O��8R�I(��=^�_�BT���K>MV]�<T�C���� ��9��!99�;6*Q�����
Q��-�������W�=�t��8͔�q�<�f�/�V(Қ]՜"sSeu��Lv�b�HHؼ�ngj�.E��Y~i�ӭ��9�F����.�n���e-��#ް��	�"��s�њ&'�z������>�+����X��j��|�@0){J�̑�F�y���p̨���k��A��HU�]!6N�'"��Rؿ�y���"N�r�?MW�:��[��턗��]�v���Mۏ+6�l�2��Y�"��2]��HqM.>.]Q��69:����)4Ƅ��u��G&4ҥ
�yLxo݆vj�8���)[{7�����AG�{�H!{u�T����aH��rw�n�W
��B|�bR$��2�u���
�e�0����PQ�5�/AQ�S3v÷�ʯ�ƚ�@u:�z�z����"W�����r�g��KCv��2��Yb~s�nw��9II6cw^Td6�7��cOTF�Ĝ�^��25?�r��cqZ��ȱ�km�M?�o�Bm���P���1�_dJ�;�8o(%s���r����Z�S p�I���&�%��;�n0�KD��H;S�
;o(�^YQw]Ю{?� �|;�i`�?kw���������|ʐ�9�H��^�D+ƣ�F�(��u�#�ܳ��������r������cE�
�7V�پ�YR����t�R�j+��[dgsl,N�Zqg�-Ȥ�8[���v��S���n�~͑��됼�j��ǜ�gB�y|C��Gn<�~p�|��Z�-����PP@���x����,�{�ٓY!	�=T�vF5I[R��/���g�N�=�6���C��م��5YL&M9Ig�)��V�'�` �w��l�X� ��ue�\���*ܴ�g�u�X��veU�+��,M2Do�5�joT؆7*���@O(�;�	0�Ȑ�~מ��A���0\E�7>��ŝNo
�5�g���R̂������01M}H*)�U|>�2���7)��������_�����i��Ƞ���Bd4||q֟�+���qkm���N�������������A���g]&w%;b���M&��Z=پ7���l�p�:��͋�~�	���?hg�"\���X��Qojq��������8�~�����%WU�3׌��_���~!H�\T� Иɣ���� 63Ƈ���M�. ihh�p���'5X~���D�h���؁r��h��\����<�Y���Ҷ|s��Sd	X2[5l�89���F��
E�!�>�{tN���J��'���;8/��p]�Q�o�� ��p;V��<#+���1����G��;>d	�nD�
Ew]Ѐ�C�K;�Sg=���lH�;��!�������������B�?����������N��IZ����n��O�����O	Ͳg�Gm�#�\^��}�IQ(�F�����:NF)Lӟ''#��������a!�28���,0�w���Y؃Eu0�s�8ѱS$�qV��>�!�ܦ^gV��'���<�9��9�����\C_�� �=8� ��*���'���6�_���g����k� Zi���P�"�@��r
mkGAI��Օ�uq��Q�հ���$�W�w5���I%u�7�Α�ey,�b2J;R	6��99R��o�Xj��ϯ	��Sٺa
�}��P8��� ��wB�)��:P��BL�i>��D�K)6GC`e^6��FϽ�4d�M��G*����}��H� �$r�h�10�����z��1����!z*ڶI4��N��s�R!�״}S��Ӕ���*]���&I�I��8���'
s����9����]	��<�)�=NeU+���YvSasb@�b��Ǭ�>��w��e����}ʲ�d|�@��6�OOƭd�cH\B�B�<���S���5�r��6x�y�3�C R	+,���*]�-U�lݭ��\/H��Ư6l�b�B�O�G����灨��n�}�`H��_�mίl^��U��-��+� ��b�'Օ���?B�����Sd?����e��&�M��� �?]u��-A�����]��XJ��Ea�UZ�������iV'Ǉ��_e��w��'�Z����?V@�OC�;n���P����4��h�;��%�^q�_ɖp��H*&��9?A�}�	���#�v�\><Z�^M��;��1�7�;�ĮW1�	(�k䭌������S�]�Ŷ��_�;ۓ8�5D���<�M�n���T2�U���/ONR
he�4E9-�w���K�NL���h$|�|��U(����l~��D�b��6����0��<�{gf=���i�u�8���}l�9��z���_{P���8��|���Jn
�)a ��R����8���w�+:=q����@D�Z��+'��!��Fj<���`�r]31lܴ-����B/���쳞+[͎��ّ-@�w��=�S�#���2<����&��Q�;	g����D�>�L@�#UP�H����
�e����5g
D�C��o������VD�=��h�a��]_�xx�}',��ʍv�g`��$�0��|�*���vx�� v���Q��VV��p��}��n���6:��#	e\���6�J:��8~W��o��$�H�%���}����cT��惕Sc�6�����՘�D���[-t!�/�'�]�L�<��X\��&Zv,D�*�gщM��+�μ�٪��~�P���\�4z��{? ��G�<�s�W�Ŭ� �^�DhG1�
��q|�>�5�mm�+���s\o���_`[����r�;�ʺ���nf�ߗ��ngx��W���ށg"�WYw[�]*��[��X<�	/Q�W� %x+�@�0�`7E� ��(Y�բqw�k_QIcr������
kJXH����|�TC�;]���wSu�XS^VT]S�J�+�|��U����ݝ�Q�*���I�9($٦���Ab����7�����G[��:3P��N� =5f�q�I�d�n���=Sz��
�|b�X�Wk�]���s��뿡� ���;����X��P���+^i��偑������Ğ��3���$J���jd�f���{�X���c	��y�e��"��Rk� #���ޭs�s�MF�E��e�B��M��i�W�� �H�b�,�T��}+�m;;z- 9�x�~��\�����B�L4�����gɴ�~UR��$r��Γ�����q���:4uª��G�2�i���5BK%3 �6�E�3�H�Mt&HwTn�+ثS��gs{~>2����x�ZȳZ�{v�$=q�[�2��M�C9��= QNGA�DE˿���\78)�� ���8�X����no�쭈	�ƾ�~	�������E�*�p  ���a�_\�sX-b�n��(���Y���H�o�i��8�����ˊ�`#�Z}-/O����W`Ȍ��9�D�|n�8t�,h�::�o�낄��l�(8��rY�IZz�����
�N�{���Ŕ£/2�n-&8b�6�s����Bp5�G�w<�h�윬�X�<�\w b�K,��C���2�B*�(�� �#�ɳ������B�UG��g	ZZl'�;��t��Z��u��$��E�5�ݙx��@��r������F���x���v�:�O�w+j��[��p�A3�م�
Lֺ��z{s�zlp�!���[IF�dfe�LA�\�'^��h��,r�IC�<	����!Wn��;�>�����N`ӃƬ����U�C"�a����$�P/q�|������w��j����P����d�"�$.�����>�t�䂧��*���g�]a�`?n�"�RSs�S���ɡ`bX�	rD��~Ub_���5��	�n�X
5��� ���<V(���j&�v��o.�dĚ$�x��-CC1ry`?ho���������|QMCECe�{eYMMo��e��_��Z�~��ggX<]�b��J��0��^�o�^�S��Qr��R��sV{Z���Z��p7m]�0��J��\g�6�ۺ`�i��J޼Y%b�������b�~��~��c��l����Y�+��� �F���%W���@>��hE�b��0�Aa1�1�!B�b"�x�ƧaM�M!�|��5HZ��(N	�W0E����?�{���y��,�N�=���{�[����=r1��^B��HD��&�_�[�;soo0�P�
r���|^]�Z+l|��`������D������s�$DoK ��r���2��P�
�(���'#T�����gT�)��_�����&6��-o�Z��H��2|M+��-)'-���h�W�E�
3�A*��O3H8��1��.� t1r�,��Z�xU�P��	��3
�%)6��=�?`z�+3�V�To�Z���c��H���2�o��-?69�D��M����K	�
a?WH���w2c�Ԕ�b�!iݮ""��]���Q3�7��O�d9ݧR�(_��$��m��1�$�1"��m�vS��a�T��T�!�ϣ�����Z���=�'�F]�kn]��RV�q\O�j�
�i�r�o@�h��|��JeOS�+����_94O�m[$5�W�=���(�B7�ϸ�$	Nd|n����8b���U;o�opy���ӫ#�]�>�~~~pA=��+e8L��+�g��քݜ���b+��Q��l�S5����mQ�U�/����	9����!mm0���"�(�s���)�$"i�͚|m�;\�@�Y��4�i�e_���;utSDq�Ʈ��]`{�zA뺘�?�z@|���S#y�+���|����c�n=�l݈y��S��6p�d(1 ��U�D<=V%TXiM!th1�H��6|���+�*1q��=2')�Bm�8�Z鹒$E6
�霓���'�w~)�Ө�����m���7\|g�4�����d�X��F���Q�U,%h��5��]��V��}	*��7MP4[C{�DiC�0G���@Q7Y�F�����Rl�m	�#�W{4��͠�����QȠ�<�[�m���ݏ�罸�Y���v6Jz�J]��RĊ�kp'fس���L��"�4Y�*�����v1,��=�}��+"e2��#��V}j��uF�f�OH��鞺.�S4g���
H��i�*�v�=oV����Jt%���F܃��gT��yLj�����J��"Ԍ~�$0�� h5x���X ��?��ڿo�b3LL5*
��Pn4�"��Iϋ%����Q��h�{
���#7�k�n�>�Ǖ��_}�t����x
�A~�@�\_[��#(gվU�py&�&���!mod/���MZ�a88Rs1��u�>G:؊s���8d�ZB�r��a<�X >b�����D�����.Y��r����5�|6+o�{�j�/��"'���@h�:��%��Fy/U^k)K��2�y4��~G���Nu�VbjB�����g�6�KV�ݰMyz�;E�#)E��E*}>C�g�4o�ލ5�ؠ����mC����~Q}���X�D]g֧!"�.Zj
���	�Ě����w`r�a|]Z�2�
���tB&Tں[n��;���6Ҭ�6hܦPSɫ�ҹ�F���.v��������A;�������w���{8�)���cZ�:��&]͌<qA�f�Fp"CI�lP����ƺ��0��dA0�:N$���격2�ԧ���(rɊ[�H��7yx0�ڂ#���$�)gkz��#���3f���5��8 ���(�H�zfY"?�����T��ɑ��p���~��Ϝh�����&��5�����zѓa�U�}�(\���Z��j+B���ʭr�a�sZ�o*hry^ǻ��(��7ip˥n3� �D��8A=H�l�,,'�6�h���b��%�CkV�$��$8�Q+�{TԔ�x�+7��B,}̜~$#���]J��2�C���S6r���yK�m+$8H3��*�!�����3��m���˸��$���#���ٶr���Yx��M������1N�}ĝ��.�=Zޔv�q�(X����B)���o�|]-�N�>9�/�W������Pt�(�����ыZ�9�Հ��|�Ҽ��|�J?)�T?���Q_ �isYI����y���	ڀ�-�N"a�������Yo��5;|׾���?#X��s{������Of.=�4����z\�7*�����$���e̥)4���s�D��&{�xǥd$��#��Xm*к����V6���h`�xy��/#���Bs�	�0�m��Ef��u }��-���Fe��8;��9�"����;�π�]�
5�i��;�"9���cad��?X�V�L9�93�_��!�����}��c�SBn{>���N0!}4$ !����Ӳ��/���ëq2��[@9�颏[y��
�	G����vYv$逘�걊��7ctX��MK@��f"*���c	�'��1 ���Bb�����Z����?'PZ����iT,d��?S����7��FBe������q�%X��V�,1�_�����9,�Q��R&�kF��� R�T�Z�-K6����F*=on�S?��a�2���f�(�.����|�D�;�Y���!ASb��_ۀ7�q��g���$�wO��j�C��"�B���q�B��b��ם����ωG��>�	t�c�[&�ef�Z���
�����'>5`��YP.�n	-��^��Lg.����,nI�sbΒ�I�>�
һF��q������x�O{�n��B�j�|��qy>��k�$�:�%Rdh�9�B-���2QT��2�0ޘ�-&N��J��מ�ݹD�7D����}��;!&���"���FGO��O�6]GXV�����Ke��C���J:�I�~@�@E4���ۙw�l��Qj����ѷ��YÓ���W�V*�m����/�x���:-�{l����Q�a�;�����捧ɀ��K�0�h�lAQ��Ć��6�>�s9|Y�~c ��h�i|�붝�Pg�G&�-"�a8S�5��+�e��+�Zg٩���������㠱kI`3���4ʐKx�
���Z�C��C�����)�P�l�,���+���l���|��ѭ�����9����$��k�}�[�k&N��>"�	�L�tx>�uH��ߕI���K/�Yn��zpi��g�T ��"��Ο2���
>D�䝩s��b;��G�d���(_D�X(������#-�w��f��*_�o/����8�,��acP�7��*%-�Lh�6��p�W�_��p�rr�{����Eʻ�%�
9�}�S�7�-K��n�95�i>m�4ⶏ��b�l��uik��#&����:�|����GyلF#�䲿�t�K�,V�����ί�f���k�G�����L��`0\�0�q�#���g��:����jT҅�e"�G�eK��b�c���sa�N SA��l����Ŏ#�`��M\c�(���n
h�t����ڇ��]��i	kk1g��gh!���<����2�6�e�k9�������H�o��{L������d����O���_���<O�3S�q����NF�!
�������|m=�qI�eB�M�X�c��Ǚ��~��ͯ�A��.�LRVp��a�bx�������<�gțG��i����~U����4��`�.x�+)�fԀo����:b4�.�!p]�y =�\[����z���21�ff1�e�ࠩ�-N#�����=TL6�0� �� �@���bso�GJo�1|Vd~�z��
��1�=�N����l����+�������D%%���m���L}zY��6
�J���Sb�,G�p4�G�����	�\�Ǵw ���۸U��+�/��B�h�g<q�O�m�{�&�5����O-cT�'��<�Q^��4Y�~66UErkCCfT8��Y��55����3��f4E<�����rg��w.�L�?(H��%��\��`RZ�i�����1P�k7�'9V,i~����n��:Ԏ�t����V�|:S�*Fǲ:�|�������7��`#4ज-��0 ������#��&��;���w�p�Z�,��b��ܖq�����s�3���*!<�� ����݌�OZ�Q�`��c��v�Ȫ'k���B�a�G��p �-�%��<2H�W�C�6;Y osK*G���	?xV��T�L�$�<��1����9{~��5ZlzK���L�Q��D�������
��g��a�3���g�סU/���B�s�E������A�G���{�(��V��*O�TU���*m��A ��g4#5$CN�'�C�O���bec5b�y��Z��x�L���O��$����=!�>P���Ix�����&�go���t}�x�JhY0t#ޣh�F ���d)/��,{��d��g����qs��̭94�<���g�ۭ�kEM�X@��29ex��+2\���8��~���{���tT8� :>' �Y)���!�xl��)�p��pYp�����eh�>.���.�<�;5�Fl�0M���%�Hd&HGeMS����Y_��>;����N�׌�[f�Fn��>aD��
��-�D�RU�Z�|�>ߒk"G��B���ER�?^}*yKJ�ȕ��/�v��$�*b-�h�M����l��+�t��|=_m_�9���!;�M�z�ߧ7$m���G	�4��)����)���8�IQ7�s�QcN�@N�逵o�q��	b*�7�C����(�q��txa��WP�������܈���͌?�O��ޔ���'��x�9�n�?kv�$I�����)d��E���~�"�`��#��&�/�՜�(����_�n"�ĳ�O.��h,�dfĩ}�uz+}.K��o������6��,(y3�FVaRZ�Y��+Ӊ![͖ԩh��8��˧����m��z�'�.B	�)�w�k`q\����ym�����F���Q"S1��(ۊz1GLj���+�ɾƠs�,��jU��h�0͟s��=6f��説�)ܵm������Q��eE�V�o<U6��g)���a���Y���Gr�l��9^)zSu��.�H�oumFѪ^A���n�>9���S���LF,ä5���/zb�{�Ү��������%=�ہȚ���t��Eo�ҩ��L�O�Z�i������s::����Q6��<��G$Is:�-���Q��:#S��̴�z�Q'249�+�UQ'qx�A�.y�����)[
�C_�p�5���7����l�|��s��$�.��P�������}Z�
�������	���Vg�7���93G�F��^?��F�7�Y�ݝRB !<k�3�J�~ak��0<vpW�����Ѓ��=
r�nx�{[^� !!)��l�����n�uѳ�����������$����Nn�S�v��)�Aw4�KT<��X�y�e�+5p�T3��d4L,�y3��UE�Z �Ȃ3�z���K�
�u�Nr^��{r�FW�����899��W��6H��͍�������
VP���,JbFy	Y�>"B�C�Wʱ� 1�mU��xz|�Bf���;!�@@�zڛ����P`�v/E��"!_Sh�`{f3�uoj�g��g?F�ѻ:Ϸ������?Cp��Kg6#��`N:4�H����\Z��`�8��L̽L՛����`g���4(@����z�u������M��i-x�����g!����o�Z����nt���A��9�H����;<��I�6Gպd,PBm�?�[���K^O�����Q��Ⲫ��ҿ��[6�F��nB) jd=r|���QE��χa<	%Q c6�j��,	��֤j� �>+�̶�䪖 `�e��1��L�e�v���v\FPP1+��G���ȿP���O�D���_�&�Y��}w�'2t��޾*�D.���hԝ��bջ'��_?�3��2<���6>3,�NK�HCi#�)L�1���/��u-�i�¤���de�z8�`��3�T_npY����f�	��PLN��OZ�3����f���p�t<�I�69ˬ�ʑ?����ܔ/�;Q�`�$ʦ�ీ�t���Lþ�::��(��'�Y��q���@�`����JI8-��*e�.�ˢ�o�;��]o�a O��u�����gD&G8�ݐ�k�!�����=�3�Y�2(x�AL2�D���D�]UN�F%�y|���:�P1�`!2H2���z�n����/�*5�R��Y)_	%%]k��3�����^� �޼�>L��;����_�Q�G)�9��:b��iL&��u~�ƙL�q&b�����rSD%MO���>�b�e�<g}�5�"*G��L�w��Ó0F��a�`�6J��q|�_D��)�팓��n_�\�=�ʍ��]���ԴT����-�[���8�=�\�i}�S�\)v��&g4�
;�����\�ci�]��CX�^�W딡�{3��6P�����/��qP�Œ,�2�в#���2b��T�a���&yy%i���&keB퀖<�p\��܈����v�]�ϲ�YG5Q���9�)tr%o�k�y��ATS�Ay� }2(-�Ǒ*����T�NFw���}l�u����&(��z�^ӯ��m�i��,`_��c�_�C�fr2>ol+�E��X�.�0��&�"Q��G�vt��D�~��P A�����P�	p7X�]�P�s��/�l �����y�L椈�4�D,aa�Q�Do���V���)�5���`tĔN��7�l&[���rbf�x%��|P���ۭ�:�5�� ����27��$��e򔅽�G�-lPwf��J���6��@?@����ȗ��@�Q@O��8:�ǣNI���`#���`-��l{�x��>�������L�o�����r��))�$�n78�ֆ�0�"bMiJ��RB�أVi[��O�+b3#�mQVW+�������
 �qk]u���@%Y���4��y�'��#�۰���S������b���%V���v��RSAt_� b�Z*Y�Q/P`�D^��m���I�L	r�8LQ�ɨ2�kQ�	G�'�~��K8ݏ���r�d��ۛ���ť�6��Mq?����U�ͱ����39#:wG�EmAN"�u��ҷ2Q�C�U�����!�:��.>Hvh�
��	[�.���˃�Fs�{ÕbY���NK{�b�9�]tڌ^�����p��FIp�A�T�JWJA1NS�w����%��}̻����4⇀�6�h���v�{�ֻ봞�ңٛq���kXK�1ɱR��P�t����se�L�c�|3݌-r����1�h���}�>��� ������"���/JU��2��U'�����?��æ�9����z�ʲ��bߐ(l��:���0Y����fT���F7���J��4��<oV�$��.��	"V|�d�$u��'h���T���=��UZP��-�v�.�6�vD.}���AYUox5CE�Ǘ� �]�;,�3I-}vu��i��>�zT�>,�uI�b��g����q=h�߼�}ȿ0��]J�akmajsG��L�Q:#�VેDB�\y�|q��RL�3���������-L�����s@���j�%�=�����z0��qAL��	A'E�NTn穭x�kx�)W"f�TVlj�
3L
-��>�aLYӄ�L�������K��N?���=Ĳ(Z��� >�}�������т���O��j{���Mh�$V�d�d�������>'b�`W�ʢ՟D���X���C�e�XN������	t�̇$,b�
4�B��P�O}�_Y-27���{���L��X[�=!��S���/?�'�B"�t���0���u87dr�Bc*�A�X|�������˶�=��3��r�%N���<�z&��'1��/k'VX���1:S��kV��R^](N��m	�g�3Ȉaq�o"%�7��%��!��S���J�DM��uz[r{���Z^]JkО��'��.�46���'�1�
`�CdHq��YOjW`p:�X�RЀ�����:�_�t��d"k�(Qڷ�מ��m/�=�IOGD7[/�T��D`g#
\��N.mB�J��X����S%�sr�'Eu=�A�BM��>�l�\�]�QtiI���|�@&��-G���Cg���,*�Hk��fW�����e�іV�)F�՝��g����[2�9R�4I��c�J����������;~��#h.E�=�~�p|lvx|c�Ӣk��L�|��U�|,m����B-�t��EϜ�7�(�߰u8X\S)*~��āE��G����{ζ_x/oj��OM��ۜY������y&)ĥ��QQ�����G��邻e�p��`ix���3�-ܶ�1���[�ۤ��I0"53�9�f��$ ��x)��C05"�`�Q�a���ԙle3x3�`E�^�ډ����=���2�@�S�i�ˏg?)����U�4QÛ��b�cD�x�h�a�Y�!ٲ�o#s��ms�B2
�o[�"�{��ޯ�@��O"o��I��Ӣp����7���?]=2��������l��tΡ�<={nh�p���y����N��$���E���5 ���8Ƽ��Q�י��  =�{��b���W	�s��C#n�M����S�y`n�I���M�5l�ɖ��t��;7y<����|�gD�/�� ���G��74��n��6�k��Y���5��r%������\�^�/�79i���V
�y��ϙ�ΖW���_}���.��g�q��K}~�}�(s5x������T2��1���?�UBםǂAE3*�?�ON��<\8sIXC�I8��3�u�鴈X z��'?2��sao�%���"3�X2�2���?vkx����\��me�����%��<�v<ޕJ��"#����B]���{�l[����K.��ߕI$2/����60��s��k	f�Y给��{vRz-�� u?�p��$'�!��Yt{!�7�oi���Aħ�ϕZ�Wh[��f��O���Ѕ�b�λ���i�KSde�U뽱�zNG.�Ȓk`(����O6�=ٍf��ӥ�q<1Ğ�Ag$~J\ȸ���׿g���l=KǍ�������B�cɤD�!q�,/lL��"V �/��[�Mɐ���@#)AHS+�8�Ne$)�]~nu�,i\=��(��r��8[y��nY�w/럽�5D�s4/e��!��Y���(�9��=bw+��r7zz�d6w�2�@P��w/Ԅyy[~��$�)�^�	����1=��02��T�P�;]P��i�	�Xȓ$r�3b��ҭ=T��}��}[,x7q!��7ԮЇz��6��؅(SX���VN�|7<�?N��<���u���m�^���b�����o+C,�_�Eh�*�JR���ȩ�?r��rU��"=�h�a��Y�D#��z<�r���F�����k�E��J�2�E�k�G�l��H{Vo�]� �`@F]H�}_�{?.�R�~��ތ�ly}���~�d �f�B�Ĥ�}Mq^�U�T%<ϡc�[?��IOᑎ���u��E���-l��5�̱c�t�w����m�OIt��9�SP��3�<PLD�m�HK���j�R��z���b�oyM�]�ۿ퉜s�&?Tr:�-H�ۨ�uFϾ<�N�J-��Ǩ9��'����T(��h�K[���Q���d�f�ܙ�N����q���e.,ηh���.pc�ԕN��������+�S����Ks�x�{�|��{���H�|����}Z�8 ��1~�@��޲)����	����ݵ����=84n�ݡ��%X�������ϝ��|9��c���c��+I���W'[ޅT����AB�afw���S vߩ3΅�#��;���w{z�yG�eL.k��h�z� �H�n<º����횞����Tx:�17��e���r����Y��/2A߁�������F�7��=�%�++��n�u�*���0\�+:8���E*!�K������pn�l��I,����,�j������E�����4��Lx<��f�u�Z�`A��x�ŉOa�d��,�����B0��]���͌:{љS['�zQC�����n��E��䣧��t�� mV��,�́�Y�G�_�w�y�Ku5H�[�q���UǺ��L4X����֞�2�jR�˚w��ק�}=B��/(����ٗQk�}?�27�P������p�����@�h�c��
�
E�Շ����mQ���Q�c0Dn���ϕĢ�WgE
��,ލcsW}d�J�6���(
I��cԈ7�E��:���� �7��d�Rw����ᄨc�����BR��|�{�@�����Gn�v[���;��E� �yS��ƍ��\zw��N��1(��xs���	����^��߄��Bi�٣�]}#��顲�B��z��R�?�In%-��:�s�^Vg-�������<Q�"�#�ҡu'���a�h#Zq>����mV$?���C�fܤ ��떍5Թ�ݎ��~�c����O��M^L��&=x�� T"�R��z֋������]9��@S�>x�s:5Ɯ�y���|>x�ғ�5)~�
D��P����[����K�W3y�6�ʄ��fa���WM��%N�}o|��yh�,��A�;V�Ia����J��+��<��R%��Yw]{���_Z ;�\��"_Ӝ��y~�Ɲ���c`a)��=\A��p63�����Y2�_�qU�zA�����W�~�r���rq*9��Pv�)i����&O�x��b���~���-˾`��ó����V(#��j�D�ꗝ�Bg)���.M�O(�Tg�}��� %4�O֍��cC2�+Ъ"J��MEC':}X���f<<][��&I-���J�凂��c��^���P�G��4߽ڢ��4I��-)��:`?�^�Y�ج�?��[3��KH���/(�G��JD�ky��	m憴����*%=I���#�mN��Ay���C��ҴA5�R�h���H8S�
Sʸ5^o�4[d¯��O�^�o����q�hb�ʳDе��,��f�	|�/-8��V��ԁ�6p�_m��K9N�Y��<��g�`	��v���NS�Q�$��p�T�烏]/��̈��ЈZ7��W����W؏�)��_9B�eo���LI��@2�i��cy����l�Ő��M�T�chjCW�۲ "؈����Bw��̀��S�YLS��ň������0eu���lUe5qO�R3�D6(۾��Di���D�=ʪf�޽��L�	7J�n,� ��g_�C�p ��3��tq��@�W�̆�k�̀�b�t�^�����㼰S�Pj�&�=6BVkvi
�fǊI>�瀈9y_z�]�j��`=�{ `s�{��
��x˱�����b0CE��R�q�F��A�~�����q��3Z�
�R\���J��Aҩ�;M����%�v�����sap`�H��2qZ���J��.��-���h����o�/���j���d(���cg�I-E�uo�F��\���G�]�ۖG��ISP��7&?Qt�4),a,��;S]h=��v1̓�<xQ{�P�mF�P�'������$�RX�뾮]+��鄾e�3�|f}��Ұ�7�ɿ<o���J���6��#K��K�dun���D���dh�3��X}B^�ٷ�sA{$��}$��= �YW�PFi�@]���X����a���2:Z�նi��k�c�_�nSjb�eǴʛ	�f��,�Zʤ_��v	��<�w
�
�5�*گz��㺎�.�'i:T����ٟ`�!��0����h9[��Y�r��Vo�+b�A8I���
b�1�N�����#����4j�ڈ��f����-� 1���*Ɲ�R�u����¨��a�oU���
���Dx<��?f!���y<7��[�H]ˮ`B^�� o����{�
P�z;,���ӵ�pe�"���?�G�,o?~h�:��5JEj��θѦL��f��>Id����d�:�ğ(����I�Kx?ܠu�M�6Fh} 1�o���E-j�!؋��v�`7�����0���ӵ&!F�ۦ{�pPG�ƤcN
E$Ȕ�����^S�M�g�z�TJ�ϓ�D�	�Gm!�`#�?f��3T��Oѭ�>!P\2����m��ݤ�ސ_��<��KߵJ%����I��	�����<�Y���<��>�"F�� -�S�^uf؍:��R������gt�x��U.*�UoJxݖY��M3��	���[�%G�=nߨih��oC[23�Z��W�$no��"�w+�e�	���2u��MQ�bwG�rdh�h��;�kb�)B��5�,}}x����O����8~����Qf�Wj��خ�*"�?���i/'��S��� k>X�M��|�℟��t�-c��(0���`�`Pw{������z=�f��8�e����F�x�c(�G���Ŧ;W����3'y����\8��T��Ӯt��F��������LN��E��}�/Zt헼�φ^#;eч/܏�.��=~d4�������Ԑ{�XL�����Lŕ�W��M��$����y&����HЂ3BJ����|�H�tG{?��L��F��49�ca�9}m8��z:�.7����jJc��5���A��&ІZd&/Hx"�R8���}�b�5���z��kޣ9 XT��&�\>5��TF��|Gi�EA���c{8$�|�O���;e�|}�ԉ�oOбJnHY/�>�phvRX*btr1�ך�/P�Ei��g z+&� ��Qk��`�L�d?����t���n�Kc���ՙ��4��i͠-0�.����D���0]R�+�$��g��A:׳6���&�)}�
���7G�(����G�D����B�����a��\Wˌ��c���)��=�[��7���U��� ��+����!�v6�4��;���fu9�3����rk��H��)���pN��y�5���!GHʅ��,�	o��S�tS���J�����ͼ�Sޖ�&��o4(�4��?#!�*0�޶���7�4:H_�����Ϭ��T��kt,��Y;���kc�`�䃧t���G��w���*�����i��+So��ڂ!�Q��2�����HC�H�0,Q:v#c3�h�����q�Z��f/�P�e��:�XA:pzJz4+Hɩt�9\�)A2�j(��p�z3�ﺠO��40l�K�@�ߪ����ٗ�`y�lY$ŷ�[������9��`��Kz���$` ���mT��|�n�����!Qp���M��N�9�1k���~�7	��`�������3\�K���^�e[w����Q�B�8B�*k���&���i&���j��O�C('����=������T��Y/��9=��M������I�.%��3�ou��N
�YT-��	A�*x�`�	>Nxt��H�bC�̧�́�nd���9����2z7����)i]�'�m����y�/�l�V��h>/wKA.}�cȟ�M_b�vL��i$�\�L_ģ���:��ˠ�i�jhkIOx�3Mq�4�c�;V��
��B�R���>�JN`��Wإ�����r�����mS�y�� ���xF*��� ��S=l���,�+~�u"@;������rka�1
�Չ��IG<�elIղ�q��{yY�;3b���Ja�D�D�����漢Ї�}���V���_�>gtFxq����L*��7��.k��}��<���B���t�߭О�x�H�x���sC�i�t7���XYnO2-i�Vzԇ)�9��X8&X�z�>˷�6��O �C���ҝ�m[��+<~E�9����B'�#��#�Ҧ�RHESD�sh��Q9���m$�J��N)4����.�[d{���$L��x�.��צ��3�'���E��kN�%O��?n)yF�Y �I65Wr��R�(W�_ah��X��v��|����.?5��*&V�)�DL����Osb4�f3��r�����yr���䈅�S�����|���á��2� ����֓���9>��U�v���+u#�J	��&���3�za�l?4A�������Լ&ŕ�IXˠ���&����t�C�����F0~��E�_��.(��g�(�/U���F���s�!o�g�M1�VO���&��z�[ �t�	���r��!\.�1�J����;ݣ�X��͟�&�w:ۮ^]@�k�K�e�8P�V?8��`� 4��[�j�R|��#5���v���(�^)�|�D�h�rG�Fj�qq,{0鿕l�������Չ,�I6�=M�㱥�j��1ψ3X� �����*&�,�ۊdרԎ!����;�aG�{���|���@Ma�,�NUƻˉ�".�@,�?=H\��?�:����Y���|̐x��3	��E���O��f��=>�,+���CŌ�Js6G����'X�)��dZ	7iz�ܗ���)j��]Ϙ=����@��Q7Jr)w�h��4��U9�n$����K/�uoP�D+������E�e�S/ߏ���jEA�@^���K�Ƃ��Han��,��(d7̷L'oʅߡD��=M%k.'�r��%���4#w
ف�TX��<�9qnz����_��g�;S�ך�{D�0�_�9E_�o�w�r_�<V�Pt��qƲ�v׽��n����7��mO���7�Up��lή�W5�"A�TI@�������M�j�GTڣ�ng䘊�TI�a��[� \��}������β����z41O����D�v]�ѷ�f��Hp�7mi�f�����)����3os�����Ft���I._}�Qg��SR��~a���}c���q����'��6��c��/~n�˱I��p����Q���-���Ⱥ�1�]gb%��M�τ)f:�q�>��#85_O���aݕ��Ģq�C˫��D|h�νE�*���w�'�*H�zppX_jG��hQ9:]EAx(ҵ����훯�������z�.��kR�K��1�tž���G�_��^l�]�7�c�����^��c�)sv]�1�?��9�/c�8<xX�+?�p����Knf��Β%6���p?�q����J-������44g�n0*�B���uP�Di�"�Ē��=v�>r"C�O5X_�z=%��M�ݿ�i�m��lg����}d�?X��:�X:��*XZ�Dw���ܝ�>� s|��#�c��w�S]��Sg��=/��Z���,\��u���H>��}�ҿ����@KǜL�(����������\WU��@�
X/<��O�w�9�@���4��f%�>�g������*�&�]�OЮy�',�fv�S�p�i���ռ��t�n��k�g|l��{>��~O�n�0����s�@�vi��$��K�� ����P\�/�2�q���}�FA��?p�e��nm1���%_R�D�,(�@+_v�rDť°ӛY��B��$"|I7 �$���%CZ�H��s`�_yȘ1G���7cO���inW��Ck�v`d �'.)j�H�P��o�����g��{ꨍ���%��W���+L�/��Rx�^Hy�{�ɰ��7�5�qf��^�m������7,~���êų��5�%3���e*��iN_6����o��{��'��J�o�Z�O����J[�BZRg����Lj(f[fj����4n �S��5�w1n�\tS�kJP�7*L�t��E�&��rI4��.���p<u��Eڿ�ޯ<����X��=�-��#r��Ej�t���x��t�iV1������wR��{��|����a�N%H��v�6���������
�Be¨�>�����6
��} .�?n��_��
I��؟N&���{X�Q���E4�����()Ň�������խI|����ï+M��X	�B��k�������ݧ�q�+�p՛D
Cy��[u� c�jh��1�m1!Hb�+^�A�9�#"�"�1�� ��"�o=־����4`��ܘ���%�
�,�1�n1�Ђ����W���k�$E f��Le��6���.��6�>8M^�J �M5��Սn:���x��<��1�+6|1�i��g5�邸�LH�iwxr�9<���Ι�4�]ӹq҇x��8\n�8����^-=ܜ�����������	w��;(�b��%f̥��>~�l�I?dW�5C~�z��������K�Y`k
�&Jo��.�^⚱ӥ������(kw���w�v�ݠ�B(���٧����˭����/���G��Ry���?%���i���ǯ]s�q�[	{�����Hvj8\ω)]�V���:7e�!�(��1-��r�3����v"���5���Ϝ�q��{��v g2p'L���р�q/�0�8=�`��jRR�wS�q9#/\��0�zљY���ad$��9���>*l�ӈ}a����EU['P�����a@~`�ߒ�>$n�$A�E�aZ�TL5�-�����x	^�:|\�h:և�)j.Ki�x,pg!��;��46P����
LZ�ծ�?�(���Mn����>BT���S��/�^)�����R���]FP�}ı[��:�3�>1����3g����x���O�Ԭ��=�)�.�Vc�!0S'9S���¥�h�`�eX���������O+"���s�G䨩�F�]��b#$�#��f��6�0�+��@�\[���2'��=Q�k]'M���pV���7�Q��}��!D����>�p_�?yMl*r���6C���<��qɥ�ò�\z�5�l|��X�v���w�Z�J��I�( 0dئ�h�_[�^���=Y�θ��Jk��֥t3���p�Iu]�r:�8!JG-�l�����Gi�Y�u�1��H5�{��k"�DAj���
RO�3�gTb���'���_���HPj---�)82��l�O��yi�u��č�_2��%����Lb�����V�#��})�ٚ�3����?�`�ldfÒ�}Qz����FI��Y:^w��x�	�
����^:�\� 
p���D%��{�SH�WO�aG�n4���s<�xv�4aH@+��;]��Ԅ�bm'�(�4w���_!� �dϲn xu*Y��,x�b�(����o��F:��t��d�e���i6��1 �k�S��D�ٟl���w�|ߗ|���`QH�n+J)���s?"W�<���6��jб��g���1��D2�R��*�%��Q�Nl���D���u�f%f5otV�Bf@�N���?�8�>Z�t�3~�O�Q�%!��aͶ���8'�b�Fl+`��O�A��E��x�.@̗���A�.)-0S��x�ҝ1��'�j��p3e_��K�����l�&zP�p�{�(2k�8�����md6h���+������a�7���k�-]Z�	qCQ%$V�3Z��a���KiEyQ}�\ ݩ\���G�
�ﻮ Q�q>�j)����I��%��]&��?�ݽ�R9ܗ��n驨����/|� �����ck�@�K�$���Ct��\N+�]v��j��`��V�3V{��'D\���9%1�<֪�����\܍�V=AZ<������0")-�b�Z���'k�v��(�9B�R C�W���wjud`l��t���������)�Q��r�5�P33s��V�<�iP�#N�RK�8d��R����}��23����F���;��MZ%e�S�2��D��,����:�W��יZ�m�`t�2�s�[��	��_L׈��J5��&�u+��xuD�F%��\1\c:�ͳHBNM��*"� �����fW�BS�D8��e$�*#�e��^8:nYok8t}�;��t����H��O�%������������֝r�s�n��������4�J�����d1W�pG��B_�����������cc�<���	7����C%e��[	�&@�gHuQ-Sʒq��I~��cr�0@�雈2[�O)�����>x[��mUc��Ѹ.�tyK�$d�N�#��S�=�HC�􁤯U�l+��Ϭ��w�,��~vd����WnK��+D�H?��p�������]��.]9��$V�GF�@̋qK}(�h���ڽ��a�&�$c���!}���Jh�vP��pq�_�Q�c��#�.�BJU�z{�9I��/����~� R`w������3�(�v�Yi+w7M�z�^�'���?�i�֑�hOrڡ�Z�2?�GF"f��[�3ym���x�6��4����|ta�ii���.�p⧘h(�R.�P���]o T�
�bc��y��JK�T�EE~#�*an+��3�ZEwE���t�������ǔ �����  ��@��Od-���쫿��*�ƬxJ(��`�F�k=��eQW$��U���4�>R���6�V� 
	��'��Y�'���Ė6��ݼ���f���ɥ���uk���FW�$`��8�Q�+a�<yKR�6�^�b>R��sVק�Ɔ4��v+�٢Q���� vH��h�.�M�hqt3�Ȩ
C�v~>��ɩ�w�x�.j�`��u�&�(<�5cN��g����t������,���bI7"��M�]g���ύ�qe�tp�@�A�A�������M111�A"O.��Ř13��Y��� lt���b\b��Nڸdt����ʕB"��e>�R����~}�owi[j���=��ņv$�~*�ޗ���(���"�GW�RπVhIUt���� ��h�c���Y<Bw�L�_:��_PQ}߀�8ۇ�"�_���gk��kI'Z4"Yd˨)?������&���]���(�yC���	��?�����c_J6|����IkpHk�,Oᑈ�6����=�A1Wƅ�u��[�SS�p݂��C��fܿ	^0�fFF"L���T)m#:MD����g��p�G������жԧX_k1��?S\T� fxf���f�����$���0��C��}r�mv�^�8�%Lnܼ.G��N���T�V�x�C92Ǿ�W_�X~��PW�k���'ŵ辋V|9��t�o��~�qU���P�Q�I}�s�����.8�AO3�B)1B��K$AE��E(9��t�SrYn�{�e���D�AW��Gl�͌\e ��B2��Fi��I�,8Cb�ܪ��s�)�vN��� A�/��#���+#֟vZ7è�%Î��t�k��_���S�w�.L��w�W���N�|�6��Ҏ�o�-� \l��!��O��Mf�;��e��(��-�_>@)�3_�=2S�X{��*A�BeIC���l�E�G���e>�2�h�誯}�H$�vhl��n����[J��e������%%��6��@�Zc� CT1��v�zaG��Y��4���y���l �ǏiC�3�UeR����0UQ�! 1f�`������Wm�馔�(Gqu2�6�I���R�� 7RmY �Ę>�6G̨�e�)�@����`\��j%c��s?��nXm//�3�?�x�O�z?��~H��䍴'�$���@��m� �|���SQ���G�3���2Ẳ.7¾�X��D��|(���2Dsx1�к��۳��i����������S�ƌ����|F�/ng�O���'��;tn����ri�vg�bK�Rv,����R�ƥ%�V�_��G�7b��ڒ�����J^{�h����Z[�pggg�G�͒�s�G\{M4Ȭ�+�J�+a����i���h��J��mk����;E��T�Q%򙒼�������y��y�SR@⦄����(�w'��Dv>�~�Ʃ�q+c���z�g&�<z߾sV���&�)g���"s�7��l��2�@��
���#�,��������2!���]�6�^�'*�q��o����R�h��H-��f��o}�ى��ux���A:�; ���(ϙ,��f���T�&Ѯ��V�����]��y��1��g�Gr�Ŭ��IM�<b���k=5�tL������r� ��e�x��Ǒ���������{LW��"�J���(�1
!�7���Z],*s�k*��u�����o������S*GQ��R|H���D�G��\� A�1�����8�ʭsaA�qb�������Kގ��������O�0����g��v��:ìz #��V{'E����[g�O��V	�U�7�c�_EP��:~C ~�MЕ��AӸtk�W�}�.-�%=dfڔ��T����s�I�MGpXD٭���6<��/�Q�<:m�;�?�w�?���g^P�Sy���x��)��q��Vj���V^*7X��X%��2x�8�#��RǦ�G+^=_j��;>­�]s�L��:8x� �Kz=�s��$#+�6ڧP���&�����	��;�M]ο�����[�ڮW}�ǳ��GY�C���;ir���Gz�DX�3�
��cE�;��jp� q��G#G��q�D�!���iK��baYTU@~.�v�-"4�N��#���"�:w�U��e
�|}tK�ɢa��4��B��/i,�+	�N����>��(<��cß��G�9�*j�%�7�☠a�Y]0�ۧ�W(+�|"��h�"e\���%�<5ʈObGS�nFm�I"�sm���,��U� i��0=�6��;�����V�Hd��K�>�~�D�\�d��@R�M�3�0N���.��.�<�zE8�R��4�Z^��u�ςn�A��չ��2�O�-AV#�f0bf*�P�ͫɺ�Cr|:Č>�L`Q0��>�
����E�Q����].Bo*�!Ƥ���k��ҳ�C�	��u�Y7D@g�@��^�G_�t�VWH��x�M1���0��.)�R_LG�~�!�#�Ό�c�0R���^���� P������ m��Adj���WgĠ��m0,�ɬa�����-_S�p�%��
Z�T�1����ﶧ0��CQlCO��+IN�βxi�t���+#��M~W&'��t0H7h���;s�80;2�7���P�4<exh�%a�@ŉ1.�^�ӡ-��g����u�*'������4�>@��=\z
Y�i�]PJ�����%T�R�۱�an&jy��K�g�n����I��]�C���@�|�μ| ߴ8q�-��A8l[��}���x)���$	D�YI��$�����ӂȮ��~q�@�G6���ٞxX����G��gÛ�jҰ�j�0Ϯ?ZB���N�s���XekO؏���cݗ�(:}��ee5�KT���?K�{�V��^�Bx4�z{Z7��~3�B��64�s�d��3x�{�+�lCֳ��מD���a�	��N�+g��������t�.���� yA���騅��Ò��yV,˽߶�Ї�d���j_9QF ���m����152 ���T\1m�3>�\@��u�L^QL=#tN��3�E�{'��N*�x���SM ����u�����������Կ�ࣀ��}��������:d��"f��Z-�A.R�f���=���A0���&��z�}~��X(c�����6�()�v[-�k��W�{��B�Ԟ��~�p�'�T�|>���c����bj�RYC[�+K�5A�����*Ѿ#����d���B�玺��}3P��tܐi���T�Tf<��:�n3�7�[ܟ��n��ۮ7W���Q����
 ��}X�%���B�Se-.緩����C@����]/!�{��݋d���?T{��4I�>wC��P�6���Y��ɉ�f�IU��"��ֺ�5�s֊}�>��d�g���ɠ��~��L�`��]S������� ��}+���stF81�0M'Z,y�^7Y!��ͫoك���U�Vd��mg�����}����g���muh�|z�F��!K�'FG6�aFޏ���&�E��]��hY����9��&3��=�j�]?E6�0���oP�B���+ڏ�)�Uߍ�Cn3Vo�D���{�d�*�a*M��mc1`�����A�A�k��*������2�}��=P�}�s�i���pzC��,�q��֮��9���w�Uύ���Y,l��� ���V\K��R��n�)���8ЀX��`� ]%b��/^��)L[t������"��Uu���x9���WM�Fe�A8̽��uᝰ�7�!J�Վ�/��u�+ܿ;�#E)��-�w
:��CbЕ"$V��h�K�R�<�>.�7���[ݷ�)3G�ϬJ\��S���/W��� ��Ru���AjO&�}`?Vt���̦bհe[�qoR�?���1�0V� ��9�B��ތ��*)�5�n��'
M�\R�N���ee�Χ��lH��Q?s��7���1�n�����r<�u�!�A%�>�[AR�>����wT�����Y�����csN���7<�&0�;N���#7�.��A�m�ft�{�3�����?�	b���h�v�bϮ�4��#�`���;�����q52D)�>�H�D]C���`Ʋez����}�^�G�<w���_¨��{ъ���Q��W8|g�~�!Qx�U����v��q��A�dҎ�=�÷�9��֫j�{� �!絴�pI�C� 猀=�j_�*�/"�O`	oU
����X�����ݎz��z��7�/4�4'�񴌦�q~Z�mG��N���k����`����&�;�2��&|��Qmn�x��eD	�1
�)�5"o�1^He���WO$�����<U�dOC�I/�2:s������~S³M��i���6{�y�LgyD�C�b���F�ލu9k��
�y�1����F���i�)�4=���?;�qY`��y3��8S��VT�P�����[yVi��s�VN����ГR�R�o���S�;(���#� ?a���!�s�y�,�a�E�a_4�8�*�|¿KX��y�Q3�ͩ�7��h�43�ۓ2��d=��3+Bш����DWe�����|;�P6�j�-�����kvf^�|��s��G!_+e�/��F�ۻ�9��[
�gԢn�_�������a�~���~	�g�K�jS'���b)%3l������_vk��J�L�����Nr-�.�̘������@�Z� }�؂�V��Oh���sHʰ��v5�z<��;�gmU�E��G��b��u���SS��� ��|`็���j������R�p)Q��|�s;+�6O�m�X�ͳN�B��^[T�4��J)K�(���:�J���j�8JF��M��*�~g�'��X���ۄt��=�࢕�����7�B�*��AW�F��N�K:h��y$11���q��Al�T��'���?Q*�#�lX�jm�b��|h�:�PD\ègs.�J�Ԑ��]8RCn��l��@=."����~'����Sx<9�P\��	0��\{yG�JJ�޼k)"dB�#q������e��ot�rH�uZ^>!�O�}�wy)z��L(��O���&U��(N {�y��S_��KN�>���~]|w���p<G��6
	�4k!gٝ�
��:�����$M��0��T[C���D��f�^v$'$s3���|ߎ�RNu�Y��ۚ�Y�pSi��PH���O���!`���}����_x0�w�.��u��ذ�n+
�<�����#J�A@�#f�U�+�3f�t @����싨^�1�j��LM���	_�8[lL
�|t�4���E�͈�El����^����/���,��Ǫ^���Q������n��:o��^dJ�B�Y./Jh��/��e�VE-�����V48�9�(��\�% �Oe'&�Af2������3yR�΃�bP�	<��㡁*���m�<+w����BYKelq2ᷤ���	��T��oN�覰��+��%;���hV�(̋h�gx�tmv"}8%I��� 2%��$�&�T�g�~���:V<�T�����"��15�ei<�-2.��{|����`�(m5xFĸ��}�'JS��|M��cr2��P�s{�MΟլ�^s��	����B8�<�%PF�����W���_r��:>e�����@/�"b�8�~�ѡ%9��OpY��Wj~6�>�+B�r�EVEi{X�駅��XZ�}zd_�>XT�%
�$�ק]�p ��H*��(KD��f���ܣ�F����K�GL�aD������o%�<#���|��r�`\��S�,B2˒=Z�F�[���PUu�"�,���Ę2�V2��`K����Ӯ�.%�8RL��"3Pox�]qˊ�9D����C&]���T�w>PB�r�k�B, ��F��p0��������wR]w�1�Lf���5Z�xxp�]_��OW�%��^��ʤd�G���Ȅ���l2ugȒ�o��2<�\��|�Pi��#�Q��4�sX/�3Ɗ��RH��@f��;=�>��K�:��^�����f\5���!)��C֣��qJ��9�6��OPB�N�l3�����jYc��6�f��o c��QC�%
��!�6�	�����+�ۑ��9BQ`�~�{��1mF�+	/P��v��ͽ,�ewA(�����	��qY=%��(��r%#����s[M�o=hlX���'�If�J��v�.W	�(;�Eh���h�ʧ��ρ}:��^����o�Z	�K'�&'�]��M��wgh�E[������1�����j#�dr�S��V�J�bb毦%i���J��o���|C#kz�)cQyt7�����>�&�֍�/�	r&���f���3�|Yo�b����fh����m����}_�]X���<<�Gw���==^T]Z���wb�50e�,T\�!���ʃ�O�ɉ���+��+MƂ�0��������|Z'��
��=8'��������»�(��w��X�A٪vIߜ�4��I!1uO���� �\~��o�I�7@j�(�{������5�U�<��K�ߒS4���!�i I�C�
��E��8ixT=nI$4<N�q�,!p>IE�p�faڸn��t��y��S��U�-�{{U�O̬��-�h�5=�*CE��k�V-{J�e��.��rK��c��-X�(�o���O�И�j)"��D�-3h�ʐZ\��B��h��k���<�w�WY�7�λt^���j�w\�ST?�u���.�RD����k�5��Jk��vnd��1*skG2���E��99e���u�\�);�=��c�v!�o��0�>�O߽��B����=��Z��W]<ͷȟ���E�<��T>�Hnd���ֿ���z`�.s�)�x�*�SR�Acx]�j��jN��.ί�.돞��e�h�>%���7��F%ꥨ�0��q�?|����ީ���b̕�x��n9�z#0���^�%O:���K��������������:�߅����wsV����)�/�Ⱦ�X������i���j��N�H} ��)`��,{�%��d�?�8Q�c�-Lr��h���Zm-�S�׷�X�?9`uk[��������}�v��z i�����p�Et�T��=FcU�Ց�[�1���NS���▯�$6�I��Z������K�箢�
�o��C�<��#$�ӰCz��]P�]��_ಛO�b:��n�'5}���G��	J��pU��'r�+]F�F�B ���K��C�,��1>�΍���ݝ4G;�K������h\z4�:4�F�g�z������G��3�u�����y�K�L����ExBF�;kii	�Օ+Bl��7������:��PX&�ݓ��W������;��k��X~K�.Đ�=����ųd/b_����>2����b���s����H����vՍqe�T�d����O�)Aqk%��̭���8>�Z��#w�N�Zm��q,����A�ȍ�e�:��	as����ߞ�{C���fAS�������7��	F��~Z�?�,Nג=�~�=qN�:���o{!⮺ȑ�|�eN_�|*�p�f%$����F:�įN4���=S�DϚ�/����0ځ�W��09Tr�Z��ġ��X���?
j���֪�ݜ{��el�6M���'�~6>[�s�-8�`z�@���F	GO��]VJya�/\�����H�H���L��p'�I,��^��������8���a㛺+k�nc۶m�wlul�6wl����f�v�6���1����j�D�ZK�?2s%>�ˡ�	���T��,lԻHCJ(��k\��(Z��Ab���v��g��0�纑uҵyi�e����fi�� 4�	^� >��'2uA���n��
sv����i�s���_�a�`�ES�AOz4!*VJ�C=59D X %ݍ5��Ā���/%_Z��.0ij bN��=X�5�;o�}��ޘ�܉���E�D^�7�[a���6��m�4x�`���E���kW�i8[��+9ao2�#i�3U��"�E���B3�DΤ�DK�)��A�NHN� �/$nis��%SLǆ�Q4����fJҿ��\s%05:��x�\��D����C���^쏴+0�Ej�� �QPGg�̉p>�.J����iV��[���0�W���J1#0'����tԖhy �~m��#1�UQ['X�·}t���J���PJ��&W��Q>��^����n|�؄�teln��}Z֬�ϓK:}��� ?��aW�mv��F�p�~�I�w��_����C/\��� V�H~<0��.4yy�Bٲ��jC&�ߍ�����@.�Ad�QM�<�%�j)���&��Ϳ)�d�q�������������!�J~�F[�����Dy�o�N2��:8N����J>O{'�NhY��&j��Ѹ�N��N��rqA�ozL,�V�!�Ǻ��ǆ}��5EFT Y$'�_loVxsW�>��]���rP�h��q~��e6|~�(�҉3��������73�{�ӭe��7H��E�~�َ�J.+"	��f� @��QE.�B����az��@���Q�rl�4ֶ7�١E$1�` _n1����b8�)�x�'�c�BȉR*̏��GQ8v�뇮�`K����]`{�p���eK�K0��%O��_�z�?\�{g�[!��{���t��,���C�Q�o!�E�h����E����~���%������2�bAb���<fs��D�h3�be�]P�=f؆�m��Su=�#�_���{�#�7(����;±};�q<s��-���h��=���⤊�ܰ��V�P1"�KB!_�В��t��3����v�p�D�d0Nd�&���`���=�f�����Xp���$iC�ݘ���XPU��N���}W}u�?�&�F���?i�^7��	/�OD��Vu�e%�'U�5���"('ӋmwAb����� &&'Yo#p=o�,�0��B�޾�����ZM���*�]��Q�KQ��t�s�FkN"�_v��3�`�����0�t�`�0��Ɠ����,��"��!@�.����fQ�v����\I)�1���"d�z��N�; g7}�soKjE�y8FMX���T֌$�_IJ�Q�'^r��jt�A�@��?[	7��ܠ�8�e�dq�A�=/�xO���������m �v5�c��{-!��8���*�JJR���+��(}��c�A5%��W��kQA�Ҕ`R%�o���e�Ɓ�}�0�������v��S����� JS;B^�/C�>�eƲ����i���s�C��n���X>3C;�����?�مH}+*�-����[LN��:�2�Ar-�G�M���@YE%x���x� �p�z���5�/�W�D<�Ҙ�L��_�~�I�4�Tq�'I��a�"�Gʓ�R�����
)���7��;��nd:YC!���7�Q Dm�q[��۹2�+�~�����1�g�^��z��Fp�+��9�3<�D]y�f�e���"��sy
��J<���<��������PZ�	�li���æ��6 �eB6��9��7<�?}�FpYp�M�	�۽##{r��&peɤ1q[�&�a����
[L���ܽ}k�Uy���<vX�q��=1Tb������1���h�
��:�/<z�Gs"�ㅐtl����X��&&y6��	(t�P�l��;���Z���h����;���jrw�Y=���H�s�#Bh舧$,�+����)����cE��8�PMeĭ������d�*���k�T��4L�ʡ�;w$�d��!'�$��a(����E�k� /f��s����~tU���Q_u_�$��#bxs�K�h��đ<o�K�ϋڲ����������>�WV��$f�gxD��۫���uL�1��Q±��T��(�0��倆I�3�� Bd[d�:#!J�������E�g���4՛L6_ʨ��������
�Q�]y�v��)*��4t�\Y�A���$�_�H��a6x
���m�Ԭ�@���s�F��2�SҦ@Z�Ud���B�'Y-trG��n9�o���8A��v�ZڛnJ^����o��DGu(�)�_�
����3��%P����@ ���-�Ɨ����N���b}N�g8����+�s��anΣY,�H�rx	9dd�Y�x�nߪq�kc��N�pUyʑE{z�?%��:��uyr�mW��h]��7�#�[���v�� ������$t��U��>�#�B}N.�?����"ⷽ�G�r��ʃ�۞�fSy����K'��ذ�V��
�	��>���K�0��^�V�z�敻	v$��3@s����T#�{���c_��V���̻3���ܠ����3� ��K��T�E�.���ʂ$Q}nn�F2������et����{"�\ѡ#�D�P1�5���>R-�
�j�h�!3�~���8�>��	UE�/����@Z�R����9S�����.O��R,��k�]g���;�3<�}��֢�J8p�A��py�U��TO�q��r��?����d���a�o��Y?�����e)��Z|%�4oHݩ���X)��N���7�á.r��"r�U�1�`Vs������8T8!J��Ug,i�1��0�a捍�����9o�p��h,�Ll�s�yV��3l�P�Ƙ�$cr��_�|�>���jpZ��kX�	5l�����zX����q���/+�~�S��0"�T$p7���7��qQ��r�ˉ�""����[��ݺ۪�Z}j(���M�3jf�`i�c�-�Z}��T%_0@+!�+5�b<4�7<I�����������3b�(&U�DN�!H7yc�&�¹G9��Tb�v�"����[qq��p�S��v��+�G��f��I�O k3��'8RULpO���% ��Ќ���V#V�'If����<Of��w��-�K:;Ks8�p�rÐS�Z��=�IE��lCL��D����^�|s0��97uޅ����$GfEה.�kV���0�4��D�!�4(�*��]Jv��1-8��LV�.�w�ˆC�-���P�q&�*Kгc�����_���&�Lzwz������������[��#������E��B��������D�`E�l=E��+#���k�&oF�\�:�+��A�_�CѼ��j��p�"�=�s�HG��Iu����ᴥ9��V�3	��D�y�w��:���Ԥ��*-�4>.���o�H��@�)C+���)EG�P[�J��Ŷ2�����ktֱ��T��*|�B-	�:���$I��BJ
�RG�Ir=qM�}��x�Gte���+� b�.b�vSU�uu�k>�^{d:c��g�w�e*��4B A�b�52���z�!�Fq��j���?�V�+�a7���gjy��6,���U;Zp�{���;���8G���
	O�T"-��K0D��Ad0�O�B�@E�6Ei���i�H0V�u�:�i�a	�af[�&�4�/�Z~�G��?	4y8�`�u�E)8f�dQq�]糉�0
�*��f'|�r�����#~�O���+(0�NB��0��N%���0��z7  ��>bZN���P�"K�

P?��H䂳@�L� n��Ômvu�ߩߊR!�i@)����	��\V�����ua!��J0������ԁ6o�"j/nMUut�Ȧo̖d��Q�|�����\��0x e��&w�WM�`�+������рϋd8�>i\,f�K��!g�V��C^�Т�l�Nk6H�_���e�*M���cKR��U��lk�_e�V�_9�j1�cǎ�pλ�lk-���`!�H��&�X�g�ԓ���g!��`���F���؍f.R�~�6rf�tP-= �+�a�qKQů�G���_K�F���I4��n��\�-r;��'��[���o�`�w�z�x�gXT���K�m4�]|�x�7�y���Y�\H�29�T�1�d�9��L�ǖ^�|,ץtl`�p!��X�u��.7����9�X���~ـ��f�����t�Y���%0�4#�NM,���Cp|x�V��$?��5Ӓ�Y��� 3�C�7>��ܠ�$)6�����/,3|�bnP��;�Pt�E�5�h��wy=��S�Ւd���v�!v\��e�6:V\Ie�}-J���̥��D�$*�q��E�#�!�A���!��DS}R�)E��	ۖ:�y2����EY��xi�G+Md�q۵TR�O~e^���u�v"1�a���ǽb`��DyE���a��=���k![#�f�IG��<���L ��<�>F��b
����n@q�a�}��Įa�?k|��:{�/�RQF��>H�35�[�G�l:��eJD��K6��	��c���e�uJ��I�A�5���pgU�3!�("#�x��Ce�p8/˖��9}��o��ܲ�}[ed������Z�k<�J;K�ş�������V�� h���\do�΍��x q���?= �I�`Q+������늎�׃po����� ƍ�1�Cÿ3�0@����@�h��A׼S�H�a�!�1��fy�ێ"7�v��ȵp��U��YT�i���8eE%�Ro�[�3f'�خc[:I�?g\5���z�I��ϫ;Hx)���)��[�Iy�IM�b��8 ����g��[�@;�I�l��(U��������H�`�P�B�`�ێ���;�af(g���Ks�	
N��Y*'��(C�26=�~*��=|M>y$:�+Znc+bQ���"Ec2�t�z1�h��Z̛��𞌚���cB6���C�����w��<�������G[��:���rm�v���X�ռTx8���UP�g��ױ��y=�״Â��j�\�8�[��]�.c�o�p�8�n�޻�F��T�K/Z�4j[M˵���i����.�}��ZJ_(��� BK)A|٘��nmS��֥F��H��vL	[(��_�$�z�ߟU.�7gTMn�:%���w�j��91����ʒU_�GGUiJ�e&��>�Ұ邧@?�Ö1��f��;���;1|gp������w,�@궼4,�T
r��F?K���38��k��U���؎��n�C�'Q���3<<ݸ(��۷����s`�L}��M�F�v�H[pƟK��5F=��/��.S�~���)U�nc�q�r�_fP@aRme��P���T�̑dˮ�Z�$6Cyq>hum���[�an(;N�|�Ԇfg ۶w'#��}B��?����I�1����ø����] ��3���}��ȳ��wr倀A� �R�-���2��<�>�'U�I3ncBm��W��4G�	*�U��L��##������5Y����j�Yr2t��e�i%=2~4Ē%�i�������JG��] �݈,��[������~o��Hc���<6q A��,H8�	��6UG�R�kJi��~lFk�Tgy6���k+昸?-%9`���+=�>�ԓ��
!Bw�.���AЛ��qe|���X��/U�^F��e�l��7��%�lL 7(�3@s��ƶ�(-rC��u�|Hw�\���`�/�a�]���!Mܬ�T6 .��L���鮷�X�t�|g)�sB�z�+xV��>�=e�Z{|b�Ĉ�$_���*|z��Gs�c�<#�����}>ʒ#��G? �S�ɷ���rY(�k��`��wr�B�M@ �}:��$󯖔a4~>��Q��u���*�F0�(���i�qM2m��F+D.�4+:r�G[���	篺:2�O��t�N��tc�5���[}U�E !�Va���ٍv#$e�g�Udbg�2Px9q'��m�H�����<�b��JW�~m�����s�p���D`�[�]�`c���T���
��V�)���g�7�#B �wJ5��|$yNPhP�̇U;����~��|!�����(������-�٪�F�|�go�YfX�oJڃ�E��"��;��x#2K�/X�r�~�P������;)�~�j�k�[K6DZ��Yf�6�)��tV8h��(O
�h��D":�Q2�Uuu�:*�`ܭ�A��1��1��_���Tf���z`�h\&F���he/|F�B�K�Y��#��k�=1k��X��O�I���K��O3��YO���J��n���hTk�Py�H����YƁr?�\�Jr�;�Ū-ߎfU����H(xM�I؎���DѢ D��r�m��B;�O������1���`�~X:\����Rԡ�<�% Kċ��֛@!r�����.w^Ne��MN�!�$�LL����[���;�Fۧ�wO����-���Ӕ	�$Z��7u6$:[�SbS68��\
|��ٻE�Y[a}(K�����/��3P}�9+��F�15T�#��k2*^-��E�����hD��z"g���*ͥ�����Gpɺ����D{�}���\.e A�逯�PNx�ڧP2�9�2�j"��+�����Ϝ����G*�l�S@)wE�6c�}E̤�]�!���D`g���������r����i����b�E�^{c:�=G�L1Su{$�"n��{���@�`��[�v;����	w6���<��f3V�#�s�!dc�	\Qtcu��*l- KȰ��ȋ[�6�{ɥv���՞��'��ʑq�2x�Ua����_��5��V6�N�qq�~��>#T=�	���%I�/jF�'�N�ۄ��-�����nly���tGO�m@ ���z��<�O7=�5�+��Q#�tyl���m�ݡ��dx��3��*8X�	�_�D�W
�p���lGҧ��R�̼�)v�۲J�-�b�F!���R8�A�J�R����F��1�E���_�X��\�@�⅌鞖�H��&��v)p�{���%�(K�n���#���my���u�͆�u�`@&*i ��F�˻d��lç�-����Zj�������
��կ�jRf^J��!�
G��*�c)��m���=Ġ�Nf'��<�7��a�Gm&m���?���·��V
�;�V�O�A��5��Q�qX��_��t?wN*
��p���϶u1K.��z\w,3�s	�48��)qI�eҺ!E&N�-O����td ��I�L�|�#@��9�� ����)����k�D4s�^����;���Y#���ѥhf�,�A ���J5�4��l�ƶ[cg+"�?�>Z���p*f5R�z�R��$�zd��_1��
,���c�,.k�M����4�}�2^�n�rds��u� ��Q�Bb��[y�Q>ǎ������u�a��y*��a\�a�9�F�Ф�2�}Z�ؕ����Bc�W�9����E�DRQ`�8b�_��*�'�
N(ɴ<��U�VͿu˻��*ʀ���twb�f#�cCaj�c�p_��m��ʶm-�Cyz۸��H���X[�Q&��]XE<<S�zx2h�L��խ��Ό15Te�kE����r*w���p��&S�0�^^�g��V�ہf� �s~of| �B�vF�z�������lu1����|��:�7X4����s/R��~�R7B#/�h͞;���4��!$`=ڌ�Kg�R���� �,#�	G	h��ZP�J���L��g��UI��7��m����ܸ��$U-_�J*H����"�r��~����w���`�\�{�t� l��|6�'g���>�w'\��7�J���ń\ܛEC]�!D�@��^ϯ�Z��('�n�?�	?��d>��Z,���>�p�!��M����`�0@��L�'i(	��'�OC�c/d� ^4$!r_m�h�`/�ލ~.��'�q�_�$���𫐎��k-��q5g.��^'����������R���y���>z�����d� 0�x֔���z��Vg���h���&���F��lvt���W
�d-�JH9L��Y�W�(�*Q/C�ȗ{�.�!^
o��w�)=���I�5�<W�<�*�4fv�n���� mC�����`ۖ�RF�G�1�Y�z�|/n*:5�_t���]��\�M/�gu�(�FN��������=696_� ����ӡQ��{su�a���w��Go��_s�/j2C��o��i��xI�FK��w��NF~, c�!h�f��JR�o1��;��|���|�4tP��"��k��$�PR:�!5iS��h(���O�ò���ȉ����ʁ��}e$xh�p���T-4�s{�w&%�/OU	gpN�,vpiLz{&T�?8 ��~8���o�k�43�"�F�=��`���[���8p�[V��p`rZXR�r�23b�E�t&6�lݚ�^lb��z�Z��
�<� |1ߢ�(p蠌)]8:�pR�"k �8 �I9[��}�6�{�S��d�x��f-�x��gU�əFh����n�mb�$��:�	��@Jq<���DWM��6G�`&z_s�3�^����K�y^ nP �^}zt?�"��G�m�����+�%XoN��h0�	&���N��Z6�jQ��Y9�s%�z��aß��Cם��ٰ��`�$E1�F�vב�&�N?��y�9�B��8Cf�"���d=eH5k�&@%?�{�&��ܻ�	W�ȅC����>\#/,n�Y}��R�2]�w�_��kM�v�-�S�=Q"�";4�K�6/=�T5C%M��G�͇��j"��\���<�l\&
�)��Y/m�^��-|q,j�m�"H��G V��*U���
�k�@p-��5W�;�3ؒ���6���	LKpS�/�^�}|�9V	���|�T����O�\�pHbV<t�,��C7�ۥ"��鬖��Ht�����T�6�yh����D��^1��h,�^�sB�<���L�C��=�Ŷ/9;5�:l������,06�̓��4��H����O=,E* i������<��d�d}7!z2��3�y�������,\��l	OK�/ǟY">?0���ly��MI�/<R��d���|$F��	��C���U�99�gFj�5��ITp\�����˚�
C��k8k�9.(��9u�m�YS��D~V&���SJm�2E^jڥ���� X��rXC' �av�+#j� x?����c!Z�s����jvz�v��֖2����4Z�Eò��u��d���?���
��� 5:��'�Dkc���z�I��2֌+���D�i��+�n�SM�����ܹכ�:�"������K$6/�9�/�}	�s��+��u��зJ�`ü7杬�c p.�	�A��6�OEU����5'�!�R7�7�ܥ�g4�.	�A�M؊ۮ��E4y"AK�n������]8\����QR �I�-!a*��G����R���_՜��lƝ+�m��j��<�|�Xl(vvvd����l�q�M����i2D��J�IB�W5��iE�\������e��YK� �xuq�x�6�E��l���2팩=�BF�7����",���]�������6�Y�2Q���(jk/��~D��z��IU���o��<�z~�R�-I���2U�ƍ6�BEE7|�3k�!��L>&�x~��g%�a��/v�C#�������"s���Ƌ���%��/��|��k�VzD�Y��p�P�����1�*�_�7����~Pk8vW�y#:���"�$�[e��Rh��#z�n�#)�{0
�X�k���y�p���f�ܴ�����K�"Xb/��*A5;bv&��L�w.`(����K��ɳLӽ�d�۠u+����rK��R�L���={,�fZ�38Sx��I}%�L~�1*�MP�3[o�$5?�?�ıA8ى�K8rsu��Hq�fx3\�EdF�po�f!�ϵ 뵁}��\��=�'�9 ������v��ˬ1��l,���E��5mNhѲ2+��v���)��?�=x��` ��Rۃ763�6��/��4��\�w�+m��ߚ��y�+*��͡�����]��j���6�
� b�I%�}����?"�2?:XƁm�/�ޚ��x�HoU������'U�`�Rt�����s��.�������Ag��4�.�'fO�)2u>U�r�dԗ��������	��V<�W@�cF��Ηx�(�ϻ����i��)�E�IB�8x�8pp�vcw}!�d��n��L��T�J��m�Us��|�HM�*�	L+����*��w� �R����L-uC;��J�v#-=���sqvg�1��ܸ�������ў��%���c�y@�d���댏8�{�hs|S����9�ΠI���Pک~���jD�V��t�~4'�)8�L��?>�J�v�q��5��!��Vo���x]��"�C�6{�y�tKy�\�ψ��[��Ϋϊ,_9���D��G�&�]��7S��W��\٪�.7h�1\/����{��D�������?t�@�0�O��N_K��ە',���S��EUv���o���Q]�1�M�jo(�(�����]}k������eoW����6�@	���K������gJ�fM�Q�*���� �+V-F�ڦ�E����7L���V�6�A�B�.^��N��D���dA�ϴ�b��!e-��{l�W!|\%���H��ù�����Wu��ǣ]�q�K�.�m#�U���M�N�՝��^/L���<T,3k���%� ���ϩ���N� �����Z.Ϗ�+�_YT@y���zBX�{�E��BR Uq;@�BW������:�Ds���?X����R����_+m�aX�F�X^�+[W�R�ȅ^�yY���F�E�Jxo߉�u��l�a���,z	��ݷZ��Ӎ=�ccT�X#1#�Qcj'^�@��PX�M�����#�	�� !}�%M�� ����iǂf�O
Rj��p���c���jf҇)^貅�g���'%�܋�|h.F�P2�89�)����!���;-oF���K4W�n�6WD����r��o��F*U�{�^v%A����Լ�Oʽf���xm3���y��#�@9����\��n���ڎ���݄�.� *0����/I"&7���}���n�L��&*�����/��:+ s��n���s�5���o�c��}ņO�"eK-���
�qQ=�`c\~�jZ��KL�R��M��;����*���+����sn�Q#C��sQu m��<N����W��jAGKأ�e�'(�H�U������̅�D�tr���IRDI ��*-ib�s;��`~F�	�YB����=�a�<Ű�>���b�J��0f��#�S�#(�ߍ(��A@�@��2!�ޮ�礢�Wr��m[�+u�b���������2hH��f�`,��(�37�\����]lU�&%��D���3�e����I�s���Ǿ�U������� �N֞����{+Z��-X�!����S�?�p�K��g�qj�5�3�	kP���o�� �ô}����h7L��Nh`氼y��`�����w+�g�%�iD�|���ru�X�I�97�e<5f+����K2F��?[[�$v��e}x��ŗ'U�i������6�
閒P>J��{Ҕ�$n��Y�_�2��۹�cyo�	�����\n�!���{��jzy�^bj
K���N�M�J��=��&�z��� ��S�%�&�bA)fvn�a�V�㴑�-:�ۙ�g!�v��ۛ����դk�~�1���ݴ�)7sV&��0�Vo1�~��}��GK� @���D]�I	�P�<����m��rÿŰq��f���A�!dƶ�� �y87(+5��خ��#�P����Q�欯�D���?��}��}�p����T��sZJ��r�%�1���pan1)�i�$(c��#�5M�Q'z$�#e����w�Ý�/�Ϗ�<�5mm�YTA���k_���y.sP8������������l�A�9��+|3�*�ƈ�߽򻎭�n 6(9�̂��A�k��{��m��S��t-���y�&�l���J2E0q��EH �ѯ�j%�x/h����r����P�����D�� 0���������kn���B�H͕�H4��&�ͮ种^$���$�_��Μl��cgX[�������͈Q�W�@Yq���L񵺝�#K2��v����~��ޥk{�d3����bͭ4��*��ɽ��k���������^��|�0��0�?3?������V_;�[�P0G�ow
�h�����uc�B��<���k^A2d2�(H�/80C.��E���ݬ�������y�Y�XZڈ����H8�� c,�0�,����*�7�e_�~ٽ�����������+Ĭ�SLcq��4��Z��B��ʼ�2�f.�A<6��`�`��d�9v��611�q�Qޕ���b}��Axã{�;W�2���r����ٳ�K?�E]�^U�?�f֓B��	���I����`��\K>J;�M��(Z4��Rb�{��1ύ*��H��vp)���rum��mW�^������Ox���&�4x@��"���RC�篶x�Z�]��"T����wB\_U:��e�	:�כ�Ź�@�Z�ۘ�h�{���Aw�uv��֦cM�xR���vG?\�l�"/��� Zޡ'�C04�7u��f���Xo)����BCV�� U&��(��{���jل�lGeY+(�DH�MH 	�sK�ueP"�G��k�����G6���;�ֲ�������Y���)�O�R��]����&>���d��������|�����H2���Z�B1�'(b|���*o�Va�b��sB�/��>dF1��>d=���m���<� ��/��D]�|`�3y�{C�q��zv�-uP���5�.��#��\?�9/�/v����p������2��],7�Q��}�$^�q��M�[}���;	ɨ�J+�j�&�	���r�G��D��l��k�rf���+:j��XB����ӰSGԓM�45�.Lﻼ٦�C*��,�v����� 
a�MT�����oi��W���M��XQM��%,�j^r��5���Z�;��b6:p)z���fGyM������B��[h�x?4�`=ٕ�Q�}��ove{��{�C q��"�ӟȧ������sfƘ���޳H�ϗ�B�!�\��u�����S�[�^���<� ܹN�o#�7��{9+��Ov�O�J��F'7*'��+�����*�	��d����6D�N4ϒ��!"����1fF`��p��U�>ApXj��{&F������V=G;%��(`}� �4?�;�5W��Q���G>2��XTƟ=i�)p����]0BP:�\Y��o�Ã�^A����ڡ�"���r��j����V��ԋ��
6���o�8�����;+���O��[�j�{��+��u��cL����.���]>����$�T�^�UV��m���l� ).������&f`�P��>h���
�Fl�����ƈ��Ͼ{8��7(�Nt$�@k�-���A�5��-͞p��d��������ߠe����h�t2�����m ��j�)
bi��kѵ��������JOt�,� �b�����G��LD�?���ZC��5�"Ӥ0��D���I$�Z�L�R ��p�8�9-�Q��O�q�\����Ӫɞ�� �u8�Y�zZ��+���xi��>Q��z���-�u����A��6���p[랯��7�f}��5�b,�[�Ȱ�é�����U����Ӆv ��Au+���?�ЧoSĀ(��_��t~8�ȇhT8(#J���ˤ��f�(�3�� f��)I�D!�՘�?��6�52�Ff1D��5�O�����+��
�	�8�g��,����Ă��E���=��!
�,�m�$�ΗV�sY5j�6t�=GO�"��HA��VB��r,>����w6 �*~Ц/ą�����TP�t�r;����0��`��מNT���rQ��X�p�����(�
;�c���*Bny0&Q����ׯ,w�i�~��]��U;�b�9EC�{�H����'�rOQX�_�=X��'/���
�*O&�O���U�$"��Tl��q��r���=�H��DS|U��t�-����x��5�A,�C���^���q���Y�8���Kbq��6�E��1��j�;�=�uT����OM4t��� ��̡�"�,!nd�
��Q�ܽY��oC'AE��[NИ����^�{��
:.;v���0eݯ�)E�_������8x�s'�M�B�o/Nx*�Y�Y5.�E�p�����W��rkey)uؿ������� �G!��,G��%��ԡ�n�E��.�[@@����Df����t��0`����5�t?W����"ߎ��n@��fu��;��\a�`5[G��:Հ�
��=H��\R�赞#��aƠ��@����/������F�e!��}\mw�l�q��R�L��B��%/��8��T� �T�i,)�5j.���v�Ҥ�����-L㈂@2<��Ϣ���X��p={�W0���Ћ�����^J�;攓Vr����qe�`?��$�w��bJ�{�]!���30�:@S�b{�5��N�p��^�g���2�f����to�믙SNٽ�����L�OoՕ��N�MS��g^ף?F)!u�X+�?���oxL$���=�I�n#B[,\w@p�BP̖�*S17�N�VD\-��7^�ؠu������38����#&OWL�\�EV�����σ��ʲ�6���v�H�h�({�6ܑ�c�j߽k�PCt�]��Y>Wy'iZ�8��6}?T$�H?�dZ�$L�(�Verǳ�p*PB7��0�\^h�B�X���jD�NC�,1R"וu�5]e5��:���������W��q���!����ݓ:Ŵ�8���#2��E���-{=�*ض�(��b��,އ��n���E�նZU�o8�d������n��Lȯt���N�G�~�xh?�����|��x~��V��Ғ�G���D�^/~v�ĜZV%Juv��--��^H��4�M��X�dY	�
)���A�q���=�iPxw�^����1�є�K����-m�om�� ��X�d��(qe��.T�Oci+�G�f�M��Td�����uC�K5��	a�j�]�Ժ���}�u���%��>���mB#�[7��&q<
�5��'�0}��+<���o{�������9��$�1�5��}Ύ������ pI�rNyj��C ��cO	�Y�eh���aEY�F;!`����Dc������<��hb��ß��}U���#���ۙ��)3�A�ǙWN���*<����LW���!�%K����2�����Ɛ�Q�^�H��
�H�8���ϥ�~K�LR�}��b�*�}����H3�nd�U�6=	m�D�SG޻zEh	V	&�F?�Y�7��K�|
mU=o�V}m��P�~<�b��9�_���a�8@��c�5M��߸ʺ��\�P;��4B��B��2�o�q��J�ލ��%cE��$�ˊm3��q�o�u�;�մ,]Cg�[�z��5x!���Rѵ}:N��A��;~������|}����A�jv����/|0Js�	 (����I���|��D뫀�'�82�&�6[���z\�U�]�/�����M��{]_щ� դD"S�&ҏ'V'��rXo�8��
�`��0�=/W)�+t�f�ZܥDK��7o��Ɖ@>w��!kܟ�e
����qhGz�@[l�lq!�n.��Un��\�^���V�NJ�w��|1_+��`�}B�}��{w�v�L �q5ޑ~������cs����X�������x�_�s)Rj�'TI��_���:--~�х����s�f�˟�#Ȱ�*��3� qo�"��W�o"?s���p�~�Y�!�t��Ӄ�y*�dF���M�H�z?s���/���������p����Hf8���ud��#Y�l�Ȉ���dIV٣lQ�q�qQ֑u�p��^G���>���ϳ������Ck		�59I�ͩ?�͏��	֜'�	�<��wFcEQ��T��]W}��V��y�d�D��x�������J���/��3v�v�������R��r�G�2�y�jb�Dni9���jf���'zw�LD�o1�~<t���$V�C�oT{&y' �3V����΋��d�i;�=ى!x��S�(Yl@�O��ǯ4-.�r��T�+�5�?T����X��W����1��|IU��;���\F�\3����K�l,zZ��Z�vU�;�ޛK�H�r��w}4G�7b5]�w?�*���H��G#�
5�}��BF�]ܾ.[z�ʠ�rL��S�\���G}�A���qM<�7�]W�5�o:��SY��4�����z|�؀:G6Y'I�Knl(�����~��:y��*q�q��UG�Ķ���[2(S3
Ѵ��M�(K��7�i����m�[.(��+	�P��/�� �OG?�6rs�ŵ�6./K��V�д�aŹ�Յ��? **j������jyYM�'���m��95PR��gj�wG�t~������|1�+�<��{~���³��ĺ���8C ���|�gx���坙�f!�"`��/�y�8:��P�+���Jb��1��T���bȹ�O�.�y���w����zo�nmQ�W7�����3G8�)��ӈ��f��H��{K��N��Ƴd[���k��k���F������_3 ����ET�cX�������@)Ŝ��b����_>RD�ϒ�0�C���ZYO����l�{�ә�ٔ�6u���e$���<b�&�^s�Y;�飨284�@<MQKg��|��3�=��*w�p���ĭ�q��5�f}`�T2n�0<$'G�_�|p� �ݩL�?��gin�p||�s��H�W����R�ҭ��wE߃��q�L2�����,�g���y��܄٤����o�%jM�ʗ�ثpq��7���C2"\eO�1),���45sB����0�5�uzx�^2z裛n�ʫ��V�l)�n^6(6�pK5���t����C���mL9H�~����dJ��9�i~�1�Q�g:�E��.���'�iQ��Ɵ,~���"�tѦp5�%�%�9����Yi)RD��u
<^�}e��w<��(��<�=[>�=�hW��`"��3���Jp���w�a��d���5n�U������bC���$�F�D8�;'�;mԍ:��'�H�nܴA�t�z�+NEp�(��4��C�Merq�8%��F�fA�i��yQ�|�ԋ���ƚL�<.��W~��b7��R�`s����6�N��9���Q��*L8x�0a��
i$R[󥤊����2B�h����#���2m�JJs�LD�bL�-����������D���G��S�r+Pn6���Q�\))d]�%#^=�1�k>}������	s�^!R�M��LwuZ'vj!��M���(��a=�I��w�K�4��վ+�ԣ�6(����ah��/an����<Va<�Y�u栴�����Ň�h��$f������'מT����],�)֝�I��;

E�ɫ�c�;�`d�8dӗh4=����5� ��w��].O��w{�l���0�s�3#.��K��e�t�����g �"�p��	��֣g���S���SҪV��y<%S�㲛�����)8˾��ЍWX8���o�ئJ��w'w_�`�Ҋ�Τ�JO�:-�ܤZ2�H�8@�EO�}'8��B�cT�1��ii9�@Ê$趯��gN��.��J�������W���JiVvgrj��F�O��h��/��qO���u�!m�Z?��ԚNޥ�g��0�>8����K��6o������k���<�=ˮ;�W�!�c����Z�����}��ӀS�;��݊����e�X��,�U�Ƒ�FY=��eF{s'[��8�IAY������ʹ�����b��w��ů3�
ˁ} v�B���,�n�:ci��_;S�ر��Ԫs�T�8�:���=N�ÏK细�%����u��b^���2�Ĉ���_EԺCW�O@������V��kL����O('�l$���`��P�`�A�|���+O�R�g��� �".?���NF�lT��7`��S �5��2?]�Dq�Y����rJZ}9� �*Ȩ�
꼸��F�D���ɭU���>1�ں��@(5�װ���?p�-5{}Ȋ��m &t�
\	�Q
9!#`֝��u�K�%�	WGš{��_�R3��2��������B��Iɷ�:?�w�查W�3h����T���;���q~�{��p*�����*��o��j�/�HQj�"���E�ȍFF��5�T�ķ���\o
�-�AE-,��$�#Ra���v�� `Uު�(T5����Lc�̐�1������+9��xs*�zQ������$�#�kj	�k6�A�-���~G�p��v�c-���鏻UA�sH�u���rQ^\}&E:5]<mQ��+0��ȭ�:_/'�J���JG�B�ׯ�;;��r�'��~=�,J�G��-���D�V	�i��y<�>:�-)j��;kxx1�"R�y��;v�)řy˓���5� �||)�j{�z�{ԓ��{��iR�O/f�������j&�?V�Y���k��-�ZT� 0�������V:�~��w{�ACMf�sB*0�b�R�1��O���,��^3�p��/цu0g�	���k^5;����Lۈwޫ/�:Q ����ǎBձ�1��/�E���)�*(Oӓ�� �N�j+!w�l�f��Nӡc�;1)l,ط�I��C���ЎO$�N��s�p��[���N(��������;��I�3X����:mf/��!A�!�3M�P"+��������{�L�-G�|�	_$��ϸ�V9;v����&VRX�R/7��}K�⁛b��O�ʗ��kVy�bF���M�x�Y���w'v�yx/�7�ɲל=)��������~�B6��c%[�.j�V3]�]�?�]tpǭ��W7=k}���~/V.ךxV��Ũ}�� ��ϳ��w�k����������p�_���C�s�@u�R�X�/UK{���od�Pz+/��&."������y�G�4�2���&~���NM��p{|j$�� R"�}P�݄+��Q��(t�^�Q~B%�+�v����g�����S/l/ �B�s�A�_��/+�ޫL�6H�&��f�^��f�w�EސVMK-�	����������p_:��[/r4��.�֍�����ra�!@��O��L�Ƿmj�,!�ct���<���NZ�e.}�"�|��Ƥt��~6�hoxj핮N��*ɭ�4�<���d+a�2x&����UyL����ْ�W�)zh�p�6��%����߿��<Ș���g�^�c��\�N�����PW�Q`�$�t�{r��U)/���ڼ�L��,z���yJ��f��3yڬ�x+�Ib�̍�?7�+n�D�wNfׯ7��ޡ��Z���շH�XŸ@�.(��s�r�_T{b��[+��r"��?���	mr�sQB���k�z�Te�ݼI�x�c�����?|kf���������v��4f�͸�"�7}m��N��PK   �z�X?�:�.  �     jsons/user_defined.jsonEQMo�0�+S�J %�u�L��i�v�P���	
����ߗ�Xo����}E�e Ԡy�p�`��v��h�� �HFce�ejQ�uݒ�'n"(1�ɇK��G�z8�i�;dul*�V�Q%�@r�*�XR^aΡ ��B�!��~����9�w��M����v0�`�i�z��jU��YE N�Z�����P�������lp�ȳʻ�DeN	�����\�\��K͋�ʽR�'x�q�u~��N��=9�QsEn�v:qy�ݘ��,Z ul�co��`,+󜕫D:x�D���6�3�b)��d������PK
   �z�X`)�t  M�                  cirkitFile.jsonPK
   5^�X�ZD) �, /             �  images/1b210ea0-4cba-494f-997a-67bd7381b5cc.pngPK
   5^�X:u�� �� /             2> images/3d480ee1-e9cf-4ef6-9de8-5a7043d7f31b.pngPK
   �z�X?�:�.  �               � jsons/user_defined.jsonPK      <  i�   