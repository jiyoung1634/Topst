PK   �|�X�IyQ#  %^    cirkitFile.json��r#Gr�_E�ޱ�u��ܭ�VX��b�X_h&�>h�� 4j$O��e�L�lp�d@t3������H����Bv��UY����n�l��n�k��Yo7�.��]��~�Ws��^o����]}�z�������ծ���6��kKu]�Y�����˪U���E]yg�1f��x���G�!����۷�.�����/��W�n��=|����p�ӑF0K+f�F0K'f�F0K/f�F0� f���3Tȅ]:��4�Yb�B$cl'����4�YVbi�C���!b@��gj��jq�D���!by���A�	["ɅI�ʒ>�	揪(�Vm�_��*Y���RA�������ғ�_BH~���)���CD
�ED"R ��򋈕_D�!"��"")dcv� 2�Jv�3�D#T� ��
\H.6 /V: �x�J�6G�f��� I�V>�rK(1�
�WUx2���3k $@h ̈CC\������%K�K�t���|\%)��\"R�o��CD
�-Qq�HQJ{z	���ˡ��[q��r+)�q�H!����B�o�!"���<{y�l	����gq/����BnD��B����˳�8�Yy���,.)�Y\��S\1��ٝ�x�k�8D� �l�R����!"��� )�Wq�H!���f�˳�8D��gqq�H!��I���q4c�G�p�|B�������8 Ty�*�#,�YZ�v����tf��9�vP:��E/���c����.�@���vP:��űV�����tfY`�+��A�Kg�%V�����tfYa����A�K����c�/�������C��� �;,��xX?������p��;,��x�	X?������<Zq��8�|�
ٍ���g��,6-X>���E�~`��#0/L�6/X>��*��i�}��������,��xX?���}�`�b���G`>^:�l_�|�3�V�A��,_���|�r�ݏ���O$�̭��xA"X~�������B���,��x'X?������W��g������|�z���`����^�������|�Ya�'�9�3�3�yr`����	�G`>^��l��|��5�`����G`>^M�l_�|�K��/?���v?����A��v?X>�q��~�~�|��B	`����G`>.� ��~�|���`����G`>.���H�Jl_<ؾx�}����K����,����
X?�}����<*���?�|i���H/�kl_<ؾ`���uv���}����+���,����X?�}�����2���,���"X?�}����$u��� �%|��J�M5#��q�-��`���#0��v?X>�q�3�~`���#0�i��/X>�q�9�~9ؾ`��ǥ��������|\�����t�h86H[ �5Uǖ�k�}s��t���l�U��yf˺�<u6���g�r��-Ȯ�}�g>.9��q�Ǚ�����<|\�v���ʶ3׀�y��x����UWg>.�:��H����%���=^��H���Q���<���7>���WYU���Cc��?N�?����ۢl�\e�/BLa�.���f�k�r�޷O}���O:��
��#7���j��m<��+�1��z�ܧ.���o���]S����)�te�?9OYM!�M����s�t��s﫲^5�κ��^�ېUm�fu�X�ڕ���'>}��ç��_��f{��-^�{�=�A��?���>�C�o��$���"P �_(������C4��1���("P �C(�]��;ᆪ%���@C
d��#(E�"�a<
b��m�%nT$3��AL��M�䍊d��=�	�p�/�tƔ��i�De�ǯ���y;��$d]��G��.+d�eq��qT$.�X���qT$.Pc��q��H\H���6`2�"6����C$�뵰<nay���H�M�A�	�):�	�I9�,�;�8ܝ���]$,��"v1���vC��8�	��]	��<�`�qT��^⠛����qT��>� &X���8*�ar,�{XGE:�O���Nw� L�<��t�}�T�ƙ��Q�������x��qT��N� &X�<�!���T��qT�î� ����`�qT��.� &X�<��t�A���9,��"v1��x��"͟�;�	�:��EDM�!?�EQa�WC��<y����f�Ƴ��Q��j���c/�G���nR�Q`�P��k��9F��bxT�������+��Q��j���c��G���n��Q`����k�a:F��
cxT����f����J�.��5h�l�A�t)�.%ۥ㻒���a���X/Z���V�~�Кt�t|X��:L�֤����"�ձa*�&�[���;B�>�:f,�?$��S�5����Hmu,�
�I7\ǇEj�c�Th�l��|����Th�l$���VǗ���d���#1_�l����VǗ��ٜ���/S�=�q=>,R[_v���]�A����#��)3*�G��ǇEj���Th�lG���VǗ��٪���/S�=��=>,rf��/S�=��=>,R[_�Bk����a����2Z������$��tE_��+���VǗ�Кt�y|X��:�L�֤����"��y^�Bkҽ��a����2Z�nD�����#��Hmu|Y�W=H_�Bk���a�+t|�
�I7�ǇEj���ThM��=>,R[_�Bkmb��VǗ�В�y��=R[��dJK�t|���e^Ǘ�В-���VǗ�В-�>��VǗ�В-�p��VǗ���1Z�3t��˼�/S�%Z����m��e*��C˵�t���e*��C�5�t���e*��C˵�t���e*��C�5�t���e*��C˵�t�U���"�ک�r@mu|�
-��r-Cmu|�
-��rMFmu|�
-��rmImu|�
-��r�Lms_�BK:�\�SG[_�BK:�\�Te~B���Thi�̍�OT����:$ʉj�3���>3ʉ��3����=3ʉ��3���G=3ʉ
�3����<�ׁ:/�����unL�=����0g{0��Q�ʳ���|��|�UE�>4��i�lCM�r��lQ�vU�2�!��U��mn��5y_�U��	,���e!�W��}<*3_�>+�xZ]W:*c��M5A�)Q0,g��(g{oS����)��e�?9OYM!�M�����.���ե��zո:�z��Y�vmVw�5�]�x�=�2)�C��C��~�����n���}���ܙo���w��C����A��C�@��з!D�@f��@�@��0���a�!2�HB
d�Q��#D(�F�"P s�bR$.k��6,o,q�"�� ���KިH�`0L��M������`L�N�$�����`L�<nay����p�o� ��-,��"q�(,�[XGE�:E0&X��<���uq`L�<nay����8,�;XGE�0&ܝܭXw�<����`L�<�`y����`y���8*�?�1���qT$^�c��q��H��Ƅ�'��)����Q�x$�	��=,��"�;,�{XGE�u^�G?�<`y����`y<��8*�c�1�n�o��x��qT$^o c��� ��H<����9,��"�|j,��<~*������{t��f@TRa%V���k2���+���e2���+���e���+��Fߥ�k���+���q�����g�����(*�&K�!
h��
�Y&��Q��j��
�Y&k��Q��j��
�Y&��Q��j��
+�	�1:�K��thyn���J�K�v��.�1^��ThI����h��ThI�����h���ThI�����h���ThI���0�h���ThI���b�h���ThI��ה�h���ThI�����h���ThI�����<X��e*��C�k�t���e*��C�k�t�Uz"��HLǗY_fu|�
-���8mu|�
-���Z>mu|�
-���Dmu|�
-����Jmu|�
-���Qmu|�
-���ZWmu|�
-���]��I:�L��thy��:�L��thy���:�L��thy-���J���+��2��˜�/S�%Z^�����/S�%Z�1����/S�%Z������/S�%Z������/S�%Z�]����/S�%Z�������e*��C˵Dt���e*��C�5Qt���e*��C˵]t���e*��C�5jt�UZI���LǗy_�u|�
-��r� mu|�
-��r�#mu|�
-��r'mu|�
-��r-*mu|�
-��rM-m��/S�%Z�����/S�%Z�q����/S�%Z�զ���/S�%Z�9����/S�%Z�����R��2:�,������ThI��k�h���ThI��k2�h���ThI��kK�h���ThI��kd�h���2Zҡ�Z�:���2Zҡ嚥:���2Z�F;s���n����r����('�xόr����('jeόr����('�Qόr����('j>��u�΋齧6}��Om�:7��L�sԯ��c,��<++_eUQ����b�:�P���m'[��]����E�yt�eu�۬qM�Wn��vˤ(gY��U�mO���W���6�Vו�ʘ�sSM�eJ���;)��������nʨn�O�SVS�sS��x�;�ˤ(gu髲^5�κ�ǯ�oCV�]��]c�kW&^ϳL����E��x۫�n�n[��/o׻�fy}U7]�\o��]��/~���3�������|u�	�}?3�32#o�r�þڢ����S������R��hF�]�T���r ΰ��s�b=;c�qJE�0����K�I)��b�Rx!��&	�T7~�%��Ȱm���2=Ƴ���M���$��Yw�1���0��uo����u�i�������������� r�_� �E��QqT_��`����R�����
�
�F�՗� �!l�?p��{>L��� ?�0���,�
�g�W��͟�Z�]cz2�d�͎�ܮ7��;�w���������v�.^��|?�[ʺ9�0���2H%a���B
q3<R�C�a
��B�S��!��dP�J�3��E*��A�r(q3L�R�C��+iR�0�ZR@v%@z��0�9bR@�%@���0�YjRq���'�
�W��!IH�&M#t$N�/M�DV�!�X�T,��[� �v�\l�X���p r��by�r���6�ѐ��!�[��L},�p�n��2����1����9<�DS�Cr�|�g�ug� ����R,/�$}H��\���;��y�)� dj���It��!�X�1�<���"��= ��cp�X  �z��Z�˒8 ��ҫ<��{'�!�X�l+��UG2��~�d[y.�xȶ�m�1�(��m ۆt|,} �W��t8�����X���<��p �o $_y.3� d��m�1�|��ms@�Mc̟���4��;Ԅ�K& ?=MF���r&勄rb��g�I�"\<�~X>�eR%����|ќ��KJ�
��G`�8� 뗔y�/���|qX �/)�*<_,���2�ڊ���G`>�L*���A�����,�꫸x��|��)��4ڐ�		M��S��]܆�}������Є<-�!ڍ�		M�S���	��Є���^��hW&L3�OmLƫ�姌�&)���#	@{B�0!�	y�>ZC�a��W�5D�0!�	y5��5ڶ�		M�+9��m��Є�
�!�
�	
ڶX�m�h�&$4!��Ak��-`BB�GU�0�m�0-�����g(�v1�bR �"e��5ahI�.LHhB^����b���&��wh�.LHhB^��=�v1`BB��E��h&$4!/�Dk�v1`BB��H�^.*���>5mj��8����W�5D�0!�	yU1ZC����WD�5D�0!�	��O/���H�v1`B^���h&$4!��k��.LHhB� ���b���&��h�.LHhB����m[���&�h�Z�Zжţm�G�0!�	�ZZC�m��K��5D�0!�	ͣ�0�}
�0�\��.�P m[<ڶ�		M��h��m��K�5D�0!�	�ZC�m��K�5D�0!�	��ZC�m��$[zAb4LG�)+\|��h�.LHhB�х��b���&��bh�.LHhB����m[���&�n`s�m��kҡ5D�0!�	�}����hw���1���9�f��z��6�e�6����̖u�y�lV�Ϭ�Pm[�]�{\�<>��8������㓚�3�O
��<>)�:���2��㓊�3�O*��<>� :���;����� ���ts<��u��U�U}���ge嫬*�����]L(O4¤�h[��]����E�Ym�eu�۬qM�Wn����ϟt��O��Bo��Ne��geO��JGeL����<�)�K?��.8��'z`S����)�~e�?9OYM!�M�����t���We�j\�u��ط!�ڮ�ꮱƵ+�nO}������bqܺ�M�c��:�M�l�e�5QJ����2~�|\]{_t�?��XL���w.x�?]�p�v��]�w�⽳x3!��1�'����}������|��?.0����)(=�x����IS�����n�����H�C��K�g|���(�Bt������J';^�O#������ϴ����y�u��F�|N�gs���9B/��8���tQJJ�m Ԣ���PPm�8��B�����'���T6Ѯ��F�)T)��8l5�BU¶»��3	!ɮ��n �&�7��2���mRBٵl�IO���s�*��	�S>8��w��W������;®�/��+���^�w/��%w��K_�w/���p�RH_��^�ӗ��%J_*�^*җʻ������*y�>�A���#�RQ�}�*�ۤ��Z>h����.��7{�0U��~}F]UѧTm����YgV��b��y������m�$�*����l����}8����j86��S@��m�͟�={�wß~�m���~ݱg���/�z��n�|�_��\ir[Yo|�pT]_Ɩ�
W��,bd�V|�FY�*Zξɳ�36����eV�3Uu����u�����"��}�i�&Y׋�v��Q��bнY��_��}��qۮ�?nA����7���T|��~���o�7�;�z��������l+�����fh�y�}���c�ŋ�����7��o������]���]�u[*������u���u��>����9~��u��vW]��m7�� 5��"��2<lpk�U�6�����w}�*�͚�/��MM���Q�O�q���yq.Be^]����p��}�w�������/�����~>Ŀ��>��{���������������w?d����g��m�6�������\��9_�Z����ι"�SW��a.m[8j)k��g��S^�Yߛ.��&����|�t�j܇��~��b�=�<��������SF����?^׻�s���c��8�W�?e����2v��r�?>�ժ[Ml֕m���!k]��:G��=��N��nJN��r� c�Tb��'d��*�x���en}U�Շ3��Ưx�������n���������z�շ������O
�L�JG0Ur�<\�������]nպ��]�U�6���>�ʮ�þ����gVӺܔ;��.�n�nҔd�/^w?ǋݳ��_�����Ac��[V�cc=x�}Sq���k�<���%����_��/���\TѧPU��o��ؙ����vc�}'������X�k��f��i�?��>�g�m�����?���H�J��_n߬��W��_}]oڛ'���}@��_�֛���{qŐO>�c/*��Þ[�x!�Vu4'�wEB����A{S6aڀp҃�i�rDM��8�g��{t��o�L����J�Ճ'=�6<����[�{*�G��~Py{���0�
|Sg��8f��U!�]���v��0e����[��z?dޢ�$k<�F���?��ϣ��u�~����n���o������ջ�Q���������?QY��k�rq�2^��������vxI�t�mZ@8�nW���,bvs���ߧ�.����r�w^��I�b_oכ������˗/|[���~��a�t�}�3�{0�s�2��>U�.�_�u}�]�޿\��}D��	���V��Bj^�Ş���8����ţ��wF���V���g5�?�ݽ8�<������n��CJw:>�u�J�aJ�����������o�y�7|�ux����3~�Ϥt�4,��~�뎁���Ô��g��fx����r�k~sn�A���ţf�q�6>O��6�ͱ���5� x���u�PM� �>Y�)�����Ի��2�p~���<��WGӿ�g��� ��
M�b?�0���p,��1jj"7%%y��.QuƔ8'�S��L2�K��K�?�>������k�E@�<���	�z� R���Nt��H�u���75����_(~�����aϺ�;<!zД�����L���}�E7x���c�T��c��������o����w���E��Oh���h����"(�2:/�e�3ɦӷ��`�л
���^����ރ��������%���z���*��c�Hiڻ���TeHꟺ@�WT�u��A�!�1xY���!i��Oyc
��k�7�J�SG�e��81�g�u�.D<���Qt���nBDR�K̰G�G<�8��(����M����]���S��WW�����n����rY�M7�/�������m}���ͷ�����+�q׻�w��O�M�[_���[��PK   �|�XWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   5^�X�ZD) �, /   images/1b210ea0-4cba-494f-997a-67bd7381b5cc.png q@���PNG

   IHDR  �  
   ��.g   	pHYs  �  ��+  ��IDATx��Y�lYv��#"#�;ֽ��z"�dw�fۂ�z2 A@����2�7���O~���h�ـX$��,H���a��������7�ΰ������9��v��*�܅��q�}�^���V!��d�������>����Q��������T6?x_�_����R�V��Kyy�R�{'�k�����L�a%�.��s�B�_��W��H��Wr��Cy��ON�˅�r��ߓ��_'������̗R�{����Z�!��b#�v+�W+�t�k�x�\��+�ڵT�B|dy�X}��R,$+2=��;��w���G�ɓ'Ooct}+��J��V�?.��R���/ˇ~��k���|�\Tr���;���L�^���ޓw�粹���ǲz�J��{�����>~(��z�gr�h./��/_zt�s���=�uG~��??�X�r�V-ձ�C��r&z�'��{�s�59��ï�lq��#����\:�]'w".��Jz����ނ�����j��v)ݺ�9;}!�z&��<?{����~p"��y"��BZ�/
i�V�O_���Ǐ9oeYJ�e:������x�(��}�:��7��ן�-�l#�oWܬ/��X�[��D��A��>(>�>�r~�J6:��:9�{"�:�|���_��O�9��ח2{�D�~��'���R�W�S�>����;"�CY|U�B!�l�:�����v/�6��Ώ�|���^�Zx�z�~�����}?�-��?��TU%y��~������o�������v-X��C����3�yt_l6<d>��ڎ�>��NV:w��5�����=��V
���[ouݗ���-��e�{m#A?ۻ�\63���̗oIY�x�A�=�#�g���8ރ�6?����ڲ}������ʂ��Ϲ�����U�=;�Ϲ�p|f}y!���4Mõy||�y����0��o���܎O5n���h���?�:��ʃ;�2S ݜ}(�j-��3y�$t�� `��Gw�J��y:ݔy)Ǉ��� Tt3�f���!�*��	l4|D��`�"V
��ذ��]hhp���s�9���x ���-s��*P ��Eč�o8?�/	���}��CX�xN����H�2W���~��ù���"�"Վ����'��o{���������F�����5F!��C��ۀ��^� }��p%���Q��U��q�\�g��r�0x�ñ�ǝ������A&�g|#�3�{q�2��k��sN���Rx���c(8;���K��> ���(�x�[�s�ysQ1�x��^2�����Bns�����7��S�ec:g�ޛ 5/S�y�@�ӥ��lͧ��=��JM��w�?�����:��?��e���3$̦kٽ��#��S:O����L�����s8=����'r;>��޿�qy���W���=~|(��������{.^-�Eu(-�F��V��^�0��T!��s%��B�%4hz�ZFj�@�ݨ���f�%##�͚��ͥ�O �jн
���sjv������ZO iW[*l�A ��e�R���37XY�h0�{i�'k#m�\Xn	�񝖚�����P��b���w{�� 	��P�v�mUY�AB �}/�;iڍ�
��n%G}�7��h���$���ތ0 �]3,�v�J��gv��_�nV|?�-�
ez�f��R����iL��k����
�ڵ�pv��Z��M�,W��"ǿ{����ϖpL�ͩ��Ϫ��I熥����٩��tWz�-��w�ST��[����=y�����H���?<�t�O0~�3*Qi�<�W|��.ikY|�b�B�h��T>��|ʍ��������Ǥ�j�zg|�)]�Y�Q��ܿ�7�E��;Sz�͡O�h��M��l\�!�àH�fΦ����������x�
������?��_�7Y������T:�tW�^��s� 3�4.U��K7���[�"pU^fR�����n"�f� ��W`\oL*�t�����n������3Y��fk]
M!��e!����X���M���m�(p�V�-��X.� i.Cb,����`�%P�{�6��\��=8�[Uxx��J\�L:����h�{XQ�Zi�`��\��+��@��:k۵�m-��J��R����J ,g�Q5��<����p?����K�.U�9�ȅ�^�B�7��yf6?�%,|1�c6���6oi�l��X�x�_S�D��]�^WJZ��j�z<��>�֫�c� �̯@�չ��<-V��n^+�+o��q�d{]��Z���:�H)�8W2��-���a�t��J� �wH���:��ν����1 ��o&
�3e�̓#�+z�
-]ߺ�U����}�����(�3�@L�^{o�s�ֆ�s>����I�;Ql�����M�MR؆W\c�=t��x��4[��k�W�"�܎O=n���`���O���}��R���+i���Rv�r�`&�6D[�wT�������B6>�E} ����A���V��-A�Q��i:�GP ��*`�¬3�6_��������V��J��
�w�n���R��{)�*\�t�[;G^u
��M�6>,^�?#w ���c��:��<#���[��,
4�,7��C���# CI�ĥśsn�=���|X�y֪�\Jޮd���f܌�Ly��E.I`��#��~..��9_���KY�_H]�%�8���g�\r-�ş��E��U�b�	xoR\nz�����X81�efJ ��9��\�|:��<*v��ߩ¢+�n� L����^�ܦQ��t�w��p��r͌�#�-S��G�QM��d�����}o:�V����y��`"�!�A1`�f�OTvt����ĵ���G��uo�$0��{�_�����$��%DOKTp�I&#@�c���MZsܗ1���tQ!IJ�����J�����<����-�~����?��y����ɱ�n�֪
�#pjm��9]�V"��ey����%��-k	x)�����K�@:nX~@��8�� |+�nUt��P9�,�H���7H�k�*���%[`���'n�`1�m4h�d���bUi�'�MsUVkV�_���Jc/��fR�jC�+/��!x�{ \��S��\�TQ����C�U)���ʖB�7 �m�V����<x��S0hl�6Y镛�W�z���
��l.�y��]D�N���$���Bu"��q���7�/_�`2;&	%���|{(y>��7����P�=�kz,��B��u���_����8�K�7��|Uq�sؘe���F��^�d;-H�]�F�2L�����@+>M��b���|������2rCX�e�v��gVP�ɣ�ʵIP� ���"s�>=�x9����2Dn��T7?���8��x=��z��;Ƃe F��~�s��t;ּ�␾G�Y����\&�ZR�����������x?��G�����fu�['�A�5���]^����\7��z��/$S�Y̜�N����]̥�*9z�m��H1W�Wz�(�Ȃ��V���T,,}E��7�"�j��3�H	U��i�1�����HڏMb$�1�� ,0$�*�:�X'ܘ���C�S8t���j�0���Z'��E���r�<���,̃�C'�y��.ޠ@�:��mĲ��u�e��h}�h������,���/��n٢4V.��$��� c��s�4b�s������fN��b!HZY��c����R�0�k�Z]f�_�t{���9U�2�7��� <��/�lp���$4��H��5<7<%b�s�'�M�j��D��u�&��[#�A��iz�	��D?�<��N�a#�� �b�y�/z_�yBLˆp ��c�u�P|4�+����y�|�DP X]&{��kŋ�׸�1�:h0�o����I���roƥEt$Kf>=�����Y�I����U�;��^��r;���x?�q�������Z���s	땬��%��R��x� � P�*7�88�l����S�7ɋ�wrW.�/�Wj	�����B3݅��3�w�UfD��48��"�;1g�;q�p���(�I���8�4�I�
{\��� Z�!�s�k( ����gnssW{�,ܥbn|e�v�%׹+��Zt1
��r����)���,^lbHL�%��"۱�p�� � ��lq?����W>�w]vtW���kVΞ��?\Di�'{��9���WAQ�DA��P�\�ђW%��������ʘ�EQ9z=�lMw5��T�H}�5���?��fׯu�R�� ��~����g5�/�/�a�\:xY�����@x�q���z�������#/ �D� ��u=َ�[9IN�j5a����ɄY|ߏ3�uj�����'���U���T�a�v_��g�x v��fJ�������9h������~��{G��k6�jpm$4�Z$NfK9<<��公t�Vj���'�ߝ�"�y:��;^ʬ�����g��L(��_��\�wT��$?��i&ܠ[�5��.��9����rrS���})'''�!�S�C^���/G�Cc�Fw3����1��� ���g�Ϛ,���@��Zj��B�l#��HU�\�x�w��J#Je��\�G�r��0������ܨ��-�?��:���h'��ݞ��)��T �˄�1�!�R'n`(3��D��y����<LY"0G�E!օ�d��	�_��0w�8o��BK�G�2�f�rs��b���uk�s38�R�P�e��B���Gg	�:�`-�rS��G!�U����'Z�x���^�=lާ�ӂ�^Kon�)�&�����ߘ+��cϪ�<�\� ���N��ES`ٷ��:�2�'�p���wpnd������Kم��Z��ߊJH"QaE�G�k�~,@��<����|aJ��O퉀ۇh�N%�.H�k[���f��<R��m�􇘒�� M|��֫=�i�(}'��4O�}OU,�O������9���}m�����\W��"i�ѥV�
� L!� )6
�ܗ��wa�u�$��-6�
J�g;��h5@V���\�b.5	29ٮ.�8��ЇхeZ�~�Qd���ؒ��b�>�[R�Uj����l&xFݕ �N���}_h�;�gq�dy{1+V&-�HD٢H�5 �g�E�:<��L�LM�����"ݵ�|��R�md�[��,	,��6Ę��]w %����a�4z� �9�ͬ^2s�(�h�g�>2ݳJ?S���B9�g�����"����Do
 Ĭ(��C�yȂL��ٰƦ�̜	�� ��(�p1$��r�c1�&)�Ļ��-����������Z��h��x-�Z�X/~�Z��k�����W� �{�8/���#H|�Q$��%�p6<�t-��K�`��g������R��17�;0e�O�������-~|�q;q��x�죿S�ݪ�-�z<GΧ
�y9#����Th\��r��"e��S��~�*\,�Л��Í���-�]��&���s����=�!���q.���r�v��IN	�<\Z���a�n6�5�=Gf����(���!���k`�t��6jE���A�G	V�GM8=�Z1|C@����DW�4����
�hy&�H�rcd	dm^��f���s��k�rTf�Xi��%[�h�n�����R�ma�G� t̎D1]G�r����MB�8ޤ^#�:g�W�S���4��p�+����x���s"�
.غ�Wo�`����;�P�?ߴS:xޥ�E+8�;��cD`��m�Q��C̅���<"VE�ւ�[�!��S�AQj,���\Vt��u�l�L�x_~ �1�d�u��Uܫ���V��t�����ݰn��2"�k?���KIڷ�/=n��s�����?������=Y��۲�J�!���M:�-e~x,n����JZ�/�o�ݡ�i�;�~���kd�!���}�G�N�蒬�\D�X}"L�(�������t�����TU�\�P����&榍�3�"$�/��-���8i���"�
sk��٬��{D)IT�
H��%��U'.
�N��"`�2ˢ���b��`��D&\ʴ/�$����ps�����=�)�W�OcR~�D��R���	*w-���s6=�k�3��)!��I��y9P(1L0�BL�2���y���B1 �EУ�W�7%Ez����U%	q^�TIq���]���a�Qa�R]�F��j^�/yt�:?�x�4v����"�a�����ЍM�CDR��V��ᘞ�|�Ve���9�Tp�c�@dЧ��zq��&A�.1�(q �>�����M�ȝ*������T!N�;e�O~wY������9��?��o]]]|��iͥ��Z6WW$o,e����"�R���K1_�:��ڈ,zT�xuK�k��7��{�6���i\��S7�1�s�֍U��&A��5�@{���l��쳣�j�0����q�r��t��ե���[Z�ƺ�r�f1��c=�n� ��a~,e�'��,�q��+B�Ә�`�F�,M.Xn�&UK���L%���q�dd$�h��2�Xe�̘l��*��>
��-x���& I��[PB��b��8�>Vc��E�[���B�n!]�<CbJG����Ұ:@7�+}�Uj=G+��eZ틇�6y�֚��X�
i(������*/��1�=�[�ʒ�aN�4�����t�n�M�<�}�,�t'���E����q��qp���+]+��՛���+i�FK����`F�s���lO���F}!nP�$�TPA·���p�� ��,��6�g�|�7x���4�~��t\��@tj������Rfa!�����C�
�
p;cm��6)j�2�K��h�
�h~ W� |CFk��-G���!X;F��Ga~?ʑ,mh۬y=��1�$b婮�M�c����}�9��e�c���E�s�Z_2Eh��ڣ2Va��Ab�	�O��ݨ�RA�!.	#H,�������ͩ.� R���Ǻ՘K��]+�-�0VVb�I�����rbǸ���0��2Wݴ�"]�Vd��L	]��<�N���t���'`=��IGf�>����`�ǒ��ü����Q�C�*y�����
Lpo���k��#*}�r�k^����d�^�7��DW�44q�~R��V;[�)���Vu��7�c�s�]�J��4#=����2�ޯTѸ��ޘ/J�]b���۵B���4�_�z���&���]��1\��O�ۿϝ�W7 �b���O9n��s�����?����gGR*����G�5�.�Y>�yv rt$��T��n���9��܇*�rnd�.�	L�v`M�fqX����$8��*����9�GY�l�25A3�U|I,�+�@��OE3�֝U��w�V!�ɲK%��N��X�z#m���X�#Ty򋽑���fC��r����c.h�ՋlHV���y���M�yC�	�;�[
{g��u�=b`}YL�B�ET7
�$��^��N�MނQ������F7�]�g����D�>1��9s*$�`� �,^#_Ų\��EnR�2Z/���5��ݐ:��c���F�^&�"�����ąlkh��L�"=�O:nrO�]&�H!��vc��w= �K�{���1��}��~(��U,�m�2U	;i�,�E��3������ي�H�Js�]�')XC��-��y�im�)m����<�*ݩ�<��nǧ���9��_�tݷ�ɼʥ��|O�~[˝�5Ax�칥ͨ�TW�+P`e�C<-X�7J����2��XJU�Y�*��rs3��裻ld؎�zV2]��ݻ�[�?	ƴ�`F �Z	S��w5�[H�Y����+2Z��$��6^�1�յ@�Q�F4���6d���Uf��huV�>�p^�y�g�H=Z3;���\�.��p��n#֘[�3u	���f�Dj�Z��o���y{�؉�퀳g��=�ȼ��yk)&S���K���4�����d������PlqK4��kT�ye1�mI�����DK|���k�*/%� �h1hA󽹹٥����<0"��mI��ԝ�:kw�X�wA�O��s�A(,p5o��;�X�C$*AF�L�!p����s��[��o�NS]�Kٻ~Rxi�k��Ʊ_�]���;>���a��'?��:o�/Pf����|.�Z���(E�_I�j��y��90����_X��4 :�l�fL�#�@`�N�e�rΎyHet#S�*`!���OpI�C.)��5~����������
p}״	ˢ�����>�3�R��Vlr}�]lNZ��F���Z���r��ݷ���)�\
����B����P��*���\����&Vk��y��*�ql䆆)#HYY[��܊[@�o��D�f�Xo=+����L�<H��1�<����Moi1�Z��������88r!k�cn�j!�"�ϥ�f�Y�.����2m��a�sjM[��J�5�*�;�bVb��O�`���y�\��~�䑀����y�]E�� xt��e����n#(M�z�\L2Ů���&����Vx+qjgk����|(݈
\�����eb���G��"�W��OA?Y�3*^]���G�潈�����ݳs�,�/�٤#�~�*�]�,�us��?eN�1_8VKc��R̚�;z�B�ۜ����s�`x�b�]g���G~Z�"�L�h���5��l��<X{߅��Tɟ�%��&�[o�_v���0�_<��G(���.�RC�[䟗Ym)8�b�-�tS44��2�c����r%�\b�j7��J�b?��B�[�ԛ�QŘ�D��S�P&�ߥ��Κ'@a��gΆ�5k1'�)�o����ߍq�������?�� �2���[���p5W�ׄ(P�`f�MU� "��V�f�'�ܬ@&HQ�0����\�����{}���5��:V|Y��sJ�ق�t�t�5�c߼��nA�x�j�G��Ůi0f���M���.q �
,0���Y�c���Bj�%F���_0�%ճv�r�%��&�&��T����4��{JjJĭa���*b7��p�7xƿ������T |�|�N�,�D�I� #����݀���϶6��X2�xuт����1!�O�F\������M]����}��4B����U���ǧ����}�{������o|���x�f���M @��5t�!������QX�h7Iհ�t�1tS)GhĽ�BBx���YGل�S�p�iԘ�1ʯ`,���bC�)�b���מ9�԰c���:n_��D���07*�IzC*̞�����
h ��5��S��i2�����M&yMQ(������cz�>E{=z�_;�\4��~(ݗ�S�E-ʱ(�56���'������b���)+nQ��㓳���V�Yk����-��q�
������b���ɤB�/��x�k>��Hl���^�~��޼|�s^S��M��v�J�&�##{S��'����`t��ld�?��x�t����0��S�w���m��)����+텽XpE��?*{z�u}k�~�q����\\|���;�|v��H@As�y%�nL�zk�V�n�b�r��3+����ʭ�?���^�E�� �U�VsxWe���l�p�c��|t��՝ط9.��������1�v�Ɵ2�{�>��ػ6D��\C���P^3R6
���Q����_6�Q`��IG%��:
E���<�齄(�ܞp�cm�)9�������U��L O��t;�'K��
M	��*bp�pS\=�%�k#�=�B��>����4?%�g��#�cO�n��c�i�v�1�H"��Y��dO�����c9B��%��\����U����L����M����χ�7���O*��1�a�yZ�D_c��s�s�����t�^�CcV��9�P�Ɗa�z����'AN�붮��	����T�,�v|�q����n�����|@(]>��6
��a&m����F��s�.�Y�����\"V��@�w�Oy��Z��/�blae�c�T`$��Ʌ̈\�l5y�|s��!�j�|Okfbd�T�
��,�wр ��ɪ�nc����jbA�|L���3�{:t�qc�I��>ѱ���a�n5� ���Er��X�/���@�:�Hz7Y���4G9��`ꂟ  a��ޜޏ.�!�]��u2��KPvAdd��c�X؃���^�d]؝`�b<(�[�ɔ�˜o�� ��H��#*0��G��G�r���d��tPdT8XeIv�,2�m}��>�~�q���^���?��'��6�Z��\�nC�7������;��e��[�{�3z:��H������f��>Ĭ'�2�{S♂n���Pnǧ�����������?�ÿ}rt �
�YU�f}�#!p�{	�ޑ>su%��~[i�6,�F��`��Q�)S���B��U�B7!��T�����pE Ixi:�%�6�7�"�.�BB����v~�qͭ�Y H�æ�˛��t��
8�6vv,��k�^���t\�G��*P"��|enyƅ57�V���s���ߧ�\,@��=�����=�2XnM0̽k��Y���.y*�m=�3��5�3^w�$ w-���]�v�~�c�g/�.���������l"tnǋbϒwY�ce3;WR ���ڊ ���-�C�3�9�z�q�L�g�X�I���3v.�s�}�ݏS�d�?�ܙ�>���q�R����9�j���Λ����׷�ܹ>�sfi�V%���U]�)��������!��+�Uzߏ�v|�q���X����~���b^JUf2�+9�ZQ ����l)��6HZ�$l�v#�R摹(B�uN3����k����~Ip�C��7�Ջ�	�۩�٪���R�(}Ԡ�]+�bM��;���כ��% IqY�1�Y�nI�4,��DkS�X���,a���,(����S*z�@���]]��67�5	A{dLg���z*��{
$.r��/6s�'@�,���Ra¬(�z��b��@A��z�.1����\�!��Y�1E)�o��~L׍�O ��@�*�5ZPk8r�&�R���e5��|��v�,ΰLߘzn�O�͏D�Aaz�;v',�1�`G����{��\����A���ց�|Y�t��5�@��{�ȥ:㙑���t����H'�-�����k��}b����3^o7rp`l����-�v|�q���h��� �v^�B��Q��jzYΎX��`VK�Z���iZ+c,��:�=ja�z��*2MC^�ېVlKЅ�:1�1��1�XL.�]H�|U{�#K%����By�I�ٮ[*սM�&xj�L9b� WZ���K�hue�o�5n�5����[�\X�LyaI͖��|7/���]̄�K� �(Xu/�Af���<\L��=����T@a(̊�%�2L	Vx�$�E�2�a�%n����ט����������x�	�X���5F���Ec����N���=>���V�X�It�F0�fY�] H�1����u㓂hz֟��6}N����Rgs�	 �eV!-��p���k��]w���i|썜1-.�����@���%�1-�q㥻�����(�^^^��|���ޗ���-�~������&,������<��}Z�}�,�E��~�f?R
9��Pa����@-�b���ཚ�b��� �c�`�*�|EY�G����\�5� vG�x.�I��E,`���%�a��c<L`�Tl��x��SOީ�v�הץ�߮7����I�G�ޢ�klz+$K���Uk�T�"|[X��e����e���\бS����Z}z��]��}�����_�7l#����w��s���td1m������z~ϟ�X����%��q�<Z󇇇rzz�s����čl������/ǚ��e��q6��j}�a�M@ͼ��- ~���W]ȶ�V;�I��C�x�Y�N\�=ױw�x�np��5���T39}v_!<�si�� }o����L��C-h�A����f�wK0�0n����<��: !�v���s��G��+��bf���i6\��a}sC$a"u��.Ow1!��GO�����[�f�"l�֏\H�2[����`�'/���u�z�����S�}���p>��/��������*�혎[�������4�lkj����w@�'6��lby?����&���µ�R�k�5i��/�sf�Yޣ�F�uhśz����l�A ��d �4��"��b���֫�s�J)�]r��Ҋ0n�����9��.cU-]WPf�87�����G�f�?�.g^/�S{?�I�JW��Fw*���|Nu���o��|��7Z����Tz ���\��b -�S���9�7��[b�������غ���C@�Z"�؍�Umf�,w `�\㻬�7>�4�a���-��a��fݝww�}_�����@�us<e,"�C*��� �R�b$�ųX���\Ê]�[��7�=�T�#^B0F���P���/��9=s�'��݉'�u�]���\���� ȍ����@�:�O8X��ط���w�}���������ޒ�,��4����Re����<5�QnLG�pQ�lH�<�p�Z(a����P#�"+Y��q��>zs ��*X�ʹ�rBA�*A`��A)���U\,"`�R�2$�)ob5'c�y3��0���\V�LfX�
WT�_�Z��i��JN"���HC���a��'�*ݼ.k���&�:��7�s;F�.>���5�@%���&�L��#N�ݔͽ?�'K�����M�ki*����V�ʢ�.�s���,c�8of ��O�y� ��3�ԯ,9 ӹ�O�{��������z���z���ߦ�M�d�V��len�x��xby��PQ�?�:�Є#����	a�Mo���kt�ο�=c�!�?�`��X���.�U�K�l|���2��"�C���@����0��x��1׺��V�n&����?���O_�]��W��]�,����������xsuU���Oʫ��Le������}��_�_���_�{����Y��y����ί�}G7�Z..V�P��S��z)��R,4����j�Ϋ����c+	�����A lM��>E�
HI�)�����1'6u�E�Z0� ��{ ?��T�纋xje�.��7�|ɲm��[�슔ǎ+V�����9���iU�akno��������#��,	���c�㵍`����Y��Q��1���|Qs���5%���X۴n�5������� ���X�{�-m�4��}(��[Rb�Ìe��$��J�+���u�����1�z��~��2B���z� @)N|���m7����~�u�=�"���X��G���D�PaMפ��Ř�\m7��C��}��}��"�ey��C[No
�_/��o��㞺ؓ+/0���O;(�v0���_?^���|��>��o�����˳Ws�A�Bŀ��{ǇGrp|,GG��\����ӟ���_��W��|��-�~F������ݬ]k�BsĠk�Z�bq"\ƨ6�ca���e� ��j�V3���JZ xt3��5�QEP�d�m����y#&1^'2�{g��3�����ݬZV��˙^��<븺����V�~�����{&�v�%L@}Լi�;"��J � ���5�1�l$�Y	N+ZO��X���I(�>qg"�I����`�e�Ś/�������s�/X�up���`9�Q��r�o��n�n;�5<GoW���ļ�,(L$�`�+��c�3���=������v�YhX�,*_.�ڊ�$e��P�blt���=�����{�
~���5�����YO���b�QS,YJt�s<�&z��w��1�}�A�s�Y�>l��j1����]�Pכ���,h�YpL�{���IU���X�`�u �e�܃��Rِ�Ҏ^���q��j7������o��w���/..~����߶}���V�Fl{y������\�<y"��淢gñ���_����s��s���7s��g0�����ڦnļԅ��%�%T���=q��Z�Ř%�G��F�ٜ*� S�utp,a�$��v]n ��t��(,}���U��u�W�p)='���jZ� ��7���d*�޲=b��q�\�n���՜�e���7�Fk �0��p�2`m,a���ͦX% �7"ON�z���N��b�;�&��B���ҽH�!� 6_ ��:$���K�Cb�_�Nu��®!)5�$,�X�$tiR�*�Z���F!ZȆF�c���6z6z�Iaֽ�\�����=�9Fr������	�
b���B��6O�+ιKka���Hm,�����Ua��r`]���{�����ޛ�O�En,��,����ڒ���x��z;k|߫"���r����K����e]˽���q��{�~�^����Y���ف�O�{�kʊ��/�����|�s�.��i��0��]�O?���z�Y�w~�w�׾�<��j��Lb�3��*���+U�U!��ϟ}����������[������ɏ���S�QZ�d�.�i���]�MQZ��ꃁKZ�M�Y]��w���o)�b��n�}͘\��+�BI��rf�fY4� M�\�T���w��
hL~ڨI�X'�!�����+�ǝ���h	�x�"a��X/�=�B�3�f,��+�
C�9���rM�}��d�(�c	�7�,�&F*��y6�B0�g�88�j�[�V~3Υ��+SKdwN���Hk)g�#��a�kXD0�b�3Q�T9c���sL�B��,6����J�[��3������)cyd��Ks�g/��lt�d�&V3��
������`�U�&w�x�$�˓��|���u��t�;Z�E�f#��ZvkU^;rl�d�K��5�\���|��c�=���(���� �3������>%D���5�����LHs���p%�Wۿ���L�z�H�z򘹾���ʡ����^���s����v�B�N�Q�Լ��|x||�e�����g\��������2�.��V�a���b��낋�9�h.�
"��ق,h,\��%���n�j�Z�!V��
�3i�Z�ٚ��u����Lx���[A	�\]�ѧƍ�z��I��.9�j�BnR�x�`ta���w4�<��3�c���lm���;+~����J�ˢ�4�.�߬�tc����q����ΑZ#hq'-7>�!�OW�b����0������Va��<:��;G2/f��E]��%�����X� �	ҽ︺o�#7VѺ	���8kt"$(@�g����M^<W�s���i��(�lTAlt}p��*���Έ�S�uF��:��]@̞��X���g������D:�f3z<��
��}O�cl;)�����J�B(e6���We֯��h����A͇�Ƙ>�s�!	�I�����z&9M�T����X:g����A*� z:jc吘��@�쩄8�Ӎב���&??*=V��H��z���!�]�9�K /-]���G/ �V_/_������3y�w��q�CpU�2F|lWct��*�2�8�z��m�G����2n��������e���n�E��u^}��_?w����Y�����i~xPK���<9���_]JUߓ@�� ��
� �f��Y�ҝ��Z@��h�<XXE�0D���9PaU�wd%K}o�r���/#/�Ś����^��܏����e��B�I��R5�颷�Y���m���
�FϿޮ�������L-�/^���٩�U�Fd���U�ȣ���bG��;+�A0��7D����%�����D�@,���L�p���lVHK����J�����r���n�J7.^�C.G�w�nk���0*�Ԧ� �-��Pe6H;�)n	�-�f�y-w�:f���
�9-�����N�j1K�VbQ!���d�%�0�"V.���>ݶ�3 ^UZ1{a��{(+�S|�tz�HdFB3K�	߷��F��νZh,�󗣒��3��K���l����S-$BU�y�3X���5�eO����zlAq`����m�mQY( �k�{�H�'K�;\��i��+$zߔ:6��-5�H���3y*'��#��V�?X�bs�9V0D��E�d�8<O9V�
���ͽ��[�SP���,#,��b˚7P t�*ۂ�E�>���NO'0�ّ,�we�Ұ��.�R�<�����l�uʬ�dP����x�g\<���0e�k$�>��3�B1!����>븆*������F� '@ؿ��ҏ�@l׺W��}�r���\��A���۬;]��\��QV������?�X�u]�Q�c��������;Ϟ={���g����������O~z�4M�w���xy��?�������?�颞��ѝ�?9::z����/E~�h����T@���������<y|��՚c�e8%�nf4��t�e �����fU�ڥ{����w��RnT αq���>�X����B!��TAILxy���E��27u���5��$6׎1I�GQ��C�l���ۇ�Xg[�ut�Yk�n�|����v��	l>S�TT�g.�5\�pX�p���l6+���*��`�ѩ��s2�]l kW�Ҩp@7�P]��?��%}�V\�Q���a�,j��x����ev��T`�h�"x���Xu�X����h0_���V�r�r!6O.�T�/����w�&/(�'�77k� ����Z<�y�1]��,����X��U���ױ
X#��3ٮ�lW�Q&CJ�S�Rk���YUW��8γ��V��ޗ!���i�k��rx|�y��J�չ<X2�1�]�	~?��&E��rK��h��<a��"ѽ�����zR�ӻ�|d�%�'��o
�*�WD"���@�}2��}=�����T�f�չR�9�����sN��]��.|T�C���f�,��*B�b�ԥY��}�^�~�3�_�׼^���"8i�<�0ײo��(��4�gs�3��7�r�`�w���0���NNN�(����|
�^�q�[ȁ{U���.Pw&���W�4n�7���{����_����Y�����|�׿�����p�����]^\|.G,������Ç�o?yr��/}������o����v��o7탾i�%�fdk���c���m�T���٪�Pm/ߨ&�fx��Oi*�2Z�&��
5�2�UH�Y��C]�(0�#���[P��6m�T��)
A.���{q?�JTQ3}���r4�K�	;��li#D��s��qF#�X�)����Ft��*�=ko^�&��D�u_�g�3���e��3����N�J�YXx�j���lQD7}Nwn�Vҭ^ɺY��qA�u�Z�:0^ς���b\�LƘ,�`.g J �ؤ���t���1�B�.��]'��9DE����!6Eǋs�EJh�c�h��%��0@��e}lZ�r�do;Z�����`6� Y	VNf�c�3�d�b�A�U�ox�K��Z�=-dc��wsq����Ρ�-+�J��ɍ�:���W�)g?� �D�2N���z�5Z�%yE]o5*��6_8������X���deJU������ѵ �*x��D� ٷ�pqΦ�������.˭��=�;v^*�P�A,�˲�:�P�g�R�2�
U�@fbl\���W��4��0q����j�:�
dm)/_^J{�y��~yx,�y�����\�o��LZ^}nզ���x�1d� S!�HWp}�0�I�cw4���ŅZ�+���k
jlT�\����z������</�[��y�˓C��<���>�R/7�Q�P�P��>?}yO�k�Ea6�oW��������oȗ����w����?�3y��9�B��T9_,����{�'�`A~gu�fIB�Dl6k��TS�.`q:�l�>,��B�n�z��l���f3�a%E66h�7z՜䂂2g�H��
�Rf�%]�I��i�XP�3d�BXw�b��/a���.�,7��g+����&0�=},o�c���?�P�9���	C\���tT�������c|�����e���*2!�+�R�.��-]���
�j�����gR�� ��""��M�Bߋ�.��% �h-���-p�,����,��FP},Dw�3y�Ɔ�|�Yڸ�V�g*]8�w�e�Rk{u �����bn��Q[~.�����B8FV�3V��t.rX>�h�g)�`�D�Z@�
��
h}uT �{)W[U��L� 
7�TA'�-�C�����r鐶ӛ���Y�Txuo��:��A+\����Jf��,����Z�.Z�zd����2�u��jt�Q���K�w�7N?�x����`��a�b��T�n����<��2�
 B)�`��D��F��f���3(-�*P>��n�#��j�ry��y�f'��i��*�..������\"�G\E�S�����KNHa��`���2�>b
P g�4�Лp��TUk�����g�չܮ:�ەʱ?�����?��Ϟ���\��?x�}IZ�K�]`�#E
mG�xa]O�3=a(�S����Ν;�ч����
֙|�-�
A�����?����<<>�61A�:����_�u�ַ�Z�Z�-�Ie����֭|�W�N��F7D���r��='�'$@VY�F�>�d���J7��k��+�V5�M0�a2��ݮh� +�Y�U ��Y4��`��7���Ӎ�|9�cO]��z۬I:��&���\�U�k|�x�grx�d���ѡ<|x_�˥ԋ"��X�QJ�����n7p����h��9��Ď�a�C[F�ټ�YAk����F���T�.�3k��z��Vn���K�R�V�3�Xb2Dpѹ��*P�M^I�h��#�/��Cn�|�Ѩu�La���u�r�A%��-���ղ �ި.Wİ؆ ���xYo��O7<�՘��p�5��:0�9��1s�=�P�ݞ.P70�	� W�zɈM���p��݃�},�阳]&2 ��0���pU�p�<�t�{��c/Ȋ�y���&����>ӗ�͟����PG�;\���K�A٫О-I�c�HUR�j^�~��تeu��XP��=X�.�z^,j�ݑ{�Q�K��i������::l宜(�TT��������(�_P���g�k���K�WTb���z�#��:#ށ�公T!���&�p��\��L��ٕZ���:��i���
f^�*)]WKS���݈��e��9^�3���<���p=�������9���z����t���..X�UNE|���n�՝�V5�E0D�5�����LI���Ȱ��^���ַ8�/_���?���]��y٪ppx �AU+d�5�b�+�9��_φ���Go�7���B�p��U���Қ.��e��G?���o=|�6�|�"�����V�ri�^�
s�0�Bְ��z�D�o?6_�E�ۉ0�1ݮ[I{y)Ŧg�e�lD-�E�p�����L�P�� �k��(/"�Q�S��(Z�W�Õ��6kY�=��顥뷶4���fYoT�����Nŧn�\7�9��R�M2�-��kU���C�P��ѿ�i-�� Xo�C�0�V-M��l����Q�dw:\�}���v�W w�*l������97pj�9M|��G{�̫ ?�ׅ��g�/ղ�U���c�sF��:9�x�\����G
���[�ִPKw�X��W��T�����:��g^�xF�������x�>���c�`y](0,�zQ3���%~�k�R-���\+0��~V��R
2<��,�Q�"\��y0F,�1���WϞK��e�j��0.n�3���ϥu[��;��ܟ��Y�i�O�|���%�A,�H�m˸�wֱ����\��
`S�L�&㔬>c��������*2ꭂ�%���lG�oF��lq@��u��+���OP����U��3*/kX���N�?�����D!mo6��3�����"���%�O>ӥ>7 /b�t�K hᳫ��{��������V�ST)��:�-d�u�dW$�!ݍ�8��q�'�QWT��t�Ō��V����~Sn����\1��<��!z���6zƜkO�w	�`D|`�l�-$l͐�H��3�Db.�5��w�$��k�����CC 1Z�����G1�ö�$�.zi�G5\����~G�ݿK߶��ޕ/��^��z�+q��{��jytB�ݬg
��Z�.Xdh��\u�.��j�`�>{���.6�Z=z�d!���4��GE�~� ���Pa_���`�`S�$$�g*`50'B��f� %��&�#֌�*�l��j	�`i�dիM�˙j��EM�cI�@����K�k��2ּm�!o�Z������i�������7��9�
h��O������&E2܍ ��x�8t0!�Y�$|���_�o�*�Ҭ�n��ѳ�����\d��
3�9N?~!A����W$W��WR��Z���ՙ���]�Bt����X�0h�t�JN�η�Rm�輫����V����g���<�8�M��^��ϗ$����9?�P`\�.?:��8;Y��\�����%�y��nu��@��]�u����{�� �x����3�P`���v||O�yM�K╂��Wr���jsE�~���g	�[�0�Y�V�^1b�-\,m< �V�No�?\J?�g������x�Uӊ�FfwU��Wz���\���u�:��U���H�Q]a���~%S�d9�
�7�΂Q\��F+<�y�p�@aA!�d�a���|����F��^/,<�/�\�P$�
�{�ui�c�eq���1.��0�xqb�����Ŀ���K�֦����ʱ"�B���ʭ[齫�K`�0F��U�Uk�82GV1��|�m?�7���c
��sQ���Tx3��eH$p�3,,׽��uJ9��I�U��^\��!���V�!���÷�׾��rtrl���8W���@)�z>ȎTU�x =d�Jgx2�܎����������[��>3Chpp%S�)Ђ$Qͬ��ܕ�i �,�v�Y���{���p�`�ߑt�
��[2=4>��
��
1��@��I�j� 5�)7H��U�&T�X)K�O��� d�Z@
f�n���䳒q�m�+�6�P�h�c*k��/.����@�;�"�qkvO����GjM���5곗�r�X�B-���=��j��1:W$AA��s���r�V`V+�J7�Ďޚ4* �������g��?�Sn4� 1�stL���1��)HܻwG��,X�R��|([�^_�P>�4����]��/.i�a|�`Z�z^�S��*;��
��E�x��C}>����E�Lq>W�U�z�Q�~��=�� ��ř��s*Q��5S���K�)�
����JM�z����@�c�YG<OT�B�p�5=[��
��B���>�vh@��^��{r�U�4�1�B5��sY�ta��-��)*8_��e��`n(�>���?s�_5+�P��zSk
�8���(����k{���ȮP����b�P���Fe8�@�Q�
u���:�&��t0����B"���@���.XkE$���Դ\�zk����`���n.�v1S�X��|�k%/DL�³�,�j��"��
L-,P�R�����TC�������k�ΰ?;~�,b�1q�=��4ʂ�V9�&�B�]-#Y�(ˡ(�X��
�Ы�R�k�X�'c��Y�Ӵ�,fbd���" ��D������C�����P(���mUY���M�.��F�M�j{�O승]G�5�d����,����=W��f+��T(�,G��(��GG����"aI���Z(����a:@��ɭ:P1?����Q����],Ok5��q���q��ၬ+
��*=�l������Z���e�t����x֍��j�:��])�]����F�v-sy������B��G
|,%��r��߹j��~��rt�D�A�;���Fz��5�)�Uy�ّU�0��� 	d�����ogО-�7#���;_Q �R�`^�`.�Q�|�7$ �/aي�zI�bA��y�p�����ѫ�]x&� Ή�6�_z��?=Ν�``*x�����V7��I	dY��q3+���t���b�)����T��CxQ ��s?�)L�D.6@��g��>����������xK��rx�mk~�Rcu��V-�v��uf�tF��4n�TƖs �需��y�s�{�b�����r� �YS�?T�bqv�YD�)I�G�M�g��VcS1RZ���+�M����r�9��4�$�$*�n������To?����'�ئ����t%h��Ŕg�{J�2,d6�ք��-�]���b�Og9��7�#��X�wk�;k�i5�q,4I���ʲ!�,s�Td�)�
2X�R��������ٯT��N����(֬%��qM�-�Flp��Kz�����||��Liĺ�Po��u)�}��է&�kPl�8<�3]�d�����CX1��ˡE�V5�#�`6��-7�d�6��U��[��t��_����K�=:Q�R�3���Ժ��t���s��+���cY�w�(�yg0����8�6��7�=���Ͷ+��L|��_��1�{���>��Z�Y( �'��ά0b�jA>z�15WT((| ��L��ͽc9T�ɓGL%b~l-�h���,��RD8c��*�S�ϯܙ��@xp|"3U"hyVH�4�8��:�8+4Y�L,?؛����<Ƒ�b�4$�����2D{>���4X���B	 �Y�-��`�����t���2��*_�� ���B- �X�8Re��b0��	�T��H,�`��`�+�I�1�8 ��*<��v~��Z٤l'-C-ӗ�k�fݱ68Sk
G ���|A���d#���9<N6(0����M��x��	��,N�Z`�Vj,�#6�K1�gt6����RaJ�7�`�a��s�O��{�#�P�	V�i�����Y,�b�w�����c����#U{@���j�����9�l(�[�+�P�-����|����l�\�1m�U�����i7��~F���8��>3~'e%L�;�&K#ȱWv�IV��'��uB�k�'e4���������|A�-������γ�/dvth�1�RA�B�Z�R�d���a!j��j	\��d��/�>�_|�\^�z!��o�U[RS��㇏��[O���̲7n�2��-�+ٰzY��s�}$��tM�,\�[��6�!��V�9�l5{��:�呂|�Y� ���(L�@�`C2�_�����o(�7�ۛ���E*�3K�בR\��!��`��F�)%�L�88�W.d���FnbyC2,��b���8�~�(A��Ҏ��U�Xd@l�"��c��R;�zK�#�0Άkh(׭"�s�B	IY�̾A��0�uˣ��b����&��E�4�h=E7'b�I��w4g͇�c�P���[�2�Pyb ��͆EGR���9+\�[wx��1ň���b�
�UY��N�bg%��c�`Ƃ�9�vl����!]c�|�r���Z�G�jrg���&����tf���E�@a5��\�����3�w
t���+�d�0*u�#0����c��%9'��Y��:]T���!]�=_.K=��z�c���kZ�:^߀���c���o��`����e8��}*=?���l}Ht]g{U:�����9����zS�S^�$N�œ����\��g$���s*M�k�P� ��}�у�����|���-w�')��]Z(m÷�Ea\�/�+�W��G_�����'��r��£�O���{����R,e���w�{|pG��<��kղ��FM<U7�X���������X�fA�1�Lq���ji��e��Y�����EWg����rg��� ��v�D]G����ZSBj�g)/)?����+P��*30�n�h�ٞ�I`)N�;O��ʳJ\�I� ���"�,����X�Y�V����5�}�����0ܗ��ɀ�n��Bv@��ǜU�9�Hھ��b��@�� �=S)tp�Ȕ��' ���N,�AX�<���0�����KE�w-6+#ʪ�$2y��᥀ MSFK����c,q��"��ެB���hi��Y���)�|*K<�2��/��X'��䱿�wC.hzM�����Y�c�����1VkeGk<~��yJTvĔ�8aT�XC+,�1_o�A��m�u�_h%U�ۿ��j|�{8��ܛ�W�d�b�~ҩ{S�1ݲ0σr���s�w[^�4�rc�3M�����/<�^n6����������#�]nZ8p1�߃�]U=I(���j��ta~�����z�W���[�<^ʼ��V����&�Dr��	z $t�n*����ds�;D+)��C���?0>!�f�c�tc��)$� �Hވ��#�NMۺ�xg�/c���FI,.�+����iS��Il	 ʦ���0Ū3���w�Բ!�F���&��3�yq��F��Z(�L�{K�]��X#~,Q����m������@K��ZI]�t����V�D��su�~��K�.ZF�5�'��x/�Q�ܲo��ľ�1�^��w6�����]a7���t��,��g��2�ǷL�1�΍�K��,]j`���!�\���M��k�E�=#=��q�`�������"?*Cq	�e*��;�_N��}P�w{�`!�{�H��Hς����H�#��>���5�"f-��� �m-Z�dpL���3Q����7�}��՘���>Gky��������'!��q����[{?�O�=�Iw��+�x���H� ���W����{\����sZv���l��`�����pV��|�~���(���)\m�}���jm��i`Lv��r�D���vdE��y�(s�����\1�^����i��X<׍B�3wj�Il�w[�Z�]*f��H��y��8}.��f&���C�o�7R8�c6c\H,��ŠH����I�����Y��.K�tT@\#S����&X�<�tQHy��9Ά�?+>���jP��Χ��o�3%r7�B>*����t��pbe�)�X�b�S0���~�kVO��b�0���+���-��gfD�.2���\��E�2Ěԩ�snqq��x��1+ZE�ٲt��ND�)f���J��n�S��0?��>?�kb�8bZO�8羅���?���ܻ����u&�@�m_�7?�u�zꊑ�fYk�,av�
F�"�ke��������oO7z�ǾE��B�έ\����3L	�N�=��M`˚b��ʊj<�/����W��u_���9- ��D2�ͦ1v�x����E��:��Y#��]Bt!6
�(,v3����a�~CLDƵ��@F$��>�R�Y��,�`�A0���g�#�%ѥ���CI �O5�y�&�Y����.����P�v#�,���L��j�?/�6KO���B"d$F��~�%��n_��Sgn�$ ��l�=�!ƫl�S��"م�o�:g�٠i�	�.tn����&�S$��M$��Ɉ}��F�&挘0a�ұ�/���9 ��\�v\g_0�8�b)������E�h"X%��Hj�8�؜܃)��0�]X1�Y[ˮ��F���=lm�����r= R|�:_Jd���W{�gJ>��7Cr���,���I6�Y�!-����HBD&�- v��9}�L�q��%7��d1g.v6q�R3�{��n��*�?�޳ǲ,���<o��4UYY���ڍfDb�H$`�/�`��G�@i���D$qDΨ5~ؾ����\fV��/�7�h��Ϲ�FTvs���n!*2����s��{�m��0��ܵ�,�o4��JN]��;/�y�K�,�>��G���5y�{�"��a���c��#r�~VZk�G�yq����s�_ε�\fӅ��B�����s�ݛ�������O*��|�U��e9�8�X+�]_�nwU�Qӄ��9����e���_UB	$�(�b�5eA�5l"R�)^�e�"7$7��ؔ�L�����2tqNnV]�T�D�)��JLN�q�M�;ܸJ��Y�S�@c�tSk�Wq��V�8�$Kj���P�7WQl�h"K���yU%&(!�����������A��4�5�:���ؠ���d*��X�%��AqE'�Hm�9|�Q��K���}ii����\�_�i)���+°@yt���P 2Y���3O�^���9��T�l�,oay�2�)+�e��Ud�#Gȋzb�dR��j&�tn�4��2y����D����7�p��Ts2��r�7+�	Eg���\yV�b�Zݳ
�Ȱ-+?'>�ѿO���_X{��������ϹD��R�Ќ���ShJ�FN�m��DG�u��>v��.y+�L�+��:c�ӵ'f��K�R��Z"no�R˯"�/�q=���ٲ�%�r�_�8���Es
����d�$p����ZVzI"�rV�t�P���V�����a^�s'�ʗ�x��"M��HH41�)5�d6U���$���3��[q��V��2�*�f��8f&��؄2�l�_j�Eu���D�z�ͽ����=-;H����%��+�{�<\��LE��d�eŪ��8 ��E�`��tV�)�U\p��By�P3�Xd���QN>3a\Q�N��n9N!yw^�cYGʰė섚��/�2}���j�<�t���ܹ^�s��p��E�I�;���l��%��g��u<r�Q[�QMF
G�5�;�.�H!l�a�\�K��tZ� �����hص��D�4�y9kX��a��Uj�aq����i��L�����R���������l�)q��5���괳���ݧ^ÅK�~�̅4��C��%>�gA��@��"-���W��[��������X��\�<��������<���t��# ��~�j���UC�(%3�M]5���;��B&ʭC�Ue%�}%^!�V~峈Cˎ6���K sFX��;D�1h ��XΞz/T�����ƟC�o�*�pEקr�;�O	TDD��Xy���/4��V�2�8��n��������8�ս*���&׎?
<���W(F��yoB'���u~Ջe���h���Q��G���E����U�1�ܹ�
�^`n��������m
%[���wY9�q�����s��e�j���v�������4�\\�)x��"�Z�ε���B���Zu�����2A<�8��{�3��u�<��Q	"G��\�����;y��!��i\�\��t"Q�Bqh"�{D����h�+,��r+�Q̕�@��h���II&��ܗY��cްbRղټW��qf\�g���Țf��&ru-�����NX�M�ո��,�G�u(���Z-��3�T¸8�G��0BK�s͐䒞����� ��J\M�pn)����'ӽ���i�����hl�6�ޜ�I�|��H��#�B��psEo����a�~L�ص��ڱ�G���p�Ώ �
���_�)�>le�"-B,A� ���/���p��N�2,�&��������׳Bب��JN���M���_��:Q�<����!3}�#ɯ}��w3_o��P��{pB��y_w��1t��o�5�._K,�2Β@�M�Y*�k���X0C�	�n.�n�L��./]�gc����
�����$��KX[&Be��u�]����^��ֻ��\�/a��T�fn�:6o0�x_�/uR����zm8��d"wo���X-(�XxS4��ucno51�%_q9�&wY��-�@�NIy���z�%77�C[>i���qOzbB���U}ňq���j�Ћ��W��R�RY�_q���)G�.^G��?\N��qrn�'�5�h��ԽO�.g8hvE蔡�����
.�K�3��>��k���B��%��#�Ǳ���d��/g�0t>��O��R�c6z BG�.ϣD$�IS��)yࡆ���Mn�_�:H�*�-��*��W��e8��gD��BC�[�5��a����Ս+��,>bB��)��E_tG2�5��eew���B�_/����;/�6A\~�?=����(+�EG3�%v^*̼T+XJ
)7��Qc��F.���S+�S0���Š '���+����B+[
'F��O�:wgnY�lU�Y��u��>iY���/�����R	Lnq��g5W�`�P���8�ן��g��2�K�$+���,�٥���q�~A��Hy�����������|%�s��fd��c�O-.4����99"�b֚�D����eg��*��+ S��b=�2�m�ۘ��M51J�Z��2O��YUP�tsUQ�fa��g��m�׈��^�c��@����1�j��ԍ<�dd�����:zհ1Cp��BG��������޼���+ٳ�S�+yC^��W�X�9�8I�Eᙈ�X����$�B�_���f\�N�ȃ�-_����T_TZ2ޯ~��^臛_8�Oj*��k)Ă+��(ץ�����ೢn�+�n ���1?ϱ[ �ҸMy����E��塹�]$�@>^�-���_V����g]�zV CW�V���늵�ܮ�L]U��(�Fq��� &aT���'t��<�������
Wb��
�C~m��Vr�@/?c�X͵�n��dK�C`V�y{q�W��t���_�/�)�����g��5��������O��� �*_��������թ禐oX\c�3.�sj� ��r_֖�$Co`dK�)��GqY�b.�[�&�V��G�����9L��{2�_�t2R��.f���{�
\%ʆ�?OÃ�Q60����~�o��f�D5��f���j�^
��^��q�ڞ�Vj��>^4�Gy�^W�C�a���C��E���.�(���=|��2ғk�<�������\W_���K��7�������_4�?��7rUqe���b ������|���+�6i>�zd`�*�p)Hh�UeKC�J,�)��Tg���=���ב��~�5POF�c�~��+K�"��>��X�:O�F�c(_�+��[���F��NKs�Y��MIQ~T>���W�,TI��9fٍ5b���!.�2��e��&@j<=��ӈV2�"W���;p1u�:��)&�����)F��;UKJt����%-�x�ߵ\"��اf�ڡn[xc+�=���~.=���,�s�g��g$+�]����V�-��0
??�N�E"���s��|݈��lJ��b��Uwr.x)#f����pȊk����t9~���^��Z�h�<xv�)��{K�#�r������8Ĥ����G��@RK�(�Дˑ��v��̊nI&��/��^}��;��S/���ױ��ҵ��P�ܓe%R��k��.+?Bo����_$��ˌH�/��Ȋ�~�J��3]�C��7(
a3�p��*T|�ͅXdk'ZzP<�t�']��6��/p���6)��^�|��=QD�Xb�!Rw�̟�����di�|���J�qr��ųb�{#�.�帗I�y�Ng�`cպ�����w��C�;r
���Z��R)2WrD��iM04&-�NT���=!pe7<���S����Q_�x�U�H>?"ˋ��l�p�D��W>'�����yb�����{s��hP"�8_��5��Q�������{��z/�;o�y��J}�6�?vjc�?m�[�U-6ny�q�.b��Vp}$���ν'�{���(� ���t���%8^zŋ�_��p��Fhq�,Y�B�8�����f��2]~�J|J_]&�ؿSG<P*��"^;�K�����@r���:����Y���ֺ�����s7箬f�d���+�fG7k�-=Cn��>�i��י��R�����N��)�����)��'�H���<K�3�|vt��C��38��D����6M�"��^�Q�#�놆C<�!�N��E�x�5��C&0�R���-��+�s��ucˌSS�qa��3Nm�h��D2\�q��v���V�D��[|2�iRs���ٳ~\WK��+H���P���k�E>�6-)�R�;/�v�¸�6M�����0�͍�;O�3�umљX���eSg+?R��X\񈨙�/��>��>�3yA�Xx/�K��5X֒��������^�ݕY]]���V�����Z�ݠ�`;K�3G�0w}ο�Y>#��W�%8^zŋ��E���P��L�۪( ���!.�FTR����nR�/�	�Y�\�$���G.1�V����Ȯ	�������߿� ��2d�dW���e���6��|��JG�!��t�2��\	PQ�q�zR�l^y�������i�����sԽ�IhBͻ5	&����f�IT-�*1Z���`ȗn��|_E�&l��B��59'R��8㟫���'X�����nM9a�p�9��|C�m)ZD����S�~7-)���ҐPqfL^�ɔK��g�����}���h;ɪQ�� ͠�$O���QR��S�ΐ�x�s�穡�P�P�
G�@!���z.!�ex�����E2WÂʑ��������h^�<���w�-
ٱ�5��=ǳϾ��K8��dlE�v�xf�Z�8���C��ֹ��!�[D�
���)MDR�+����p="U��$���S~���K�]�&�˴&1�3��d�k�z=������3=0���띰�'���d"��}]^{�5'�H�����g:�^Y��YȋPV�%8^zŋ��,+���|Q|�|p3p�qE���NxV�ǜ�n@I�"a[�5�,\�U�U�f^����_��Ps���s}���)�^`����E���^��=�G�w�t�����bkAf��֖Ϻ�x_Z��b�A�mx����������m���$.;9�W�	�R�Sx��.x�,�2G�*t��2�o��;]_܇2ey��e�.p�66��o�<$R�����N��u�����?��w��Zݿ�e*�y���G�=��ACE˸[YQy�U���y�6��U-�I�B3�$ƥ��-���9<J��S�>��������,i�lY!�/��7ru��,2�i����r�.b��S�{�ZDʑ�wJ�=�p�5���l��iOC׵G�i�y;*�P9�I'�D<��1K=)��������bZ��u����E�]����j��H7dW���n�Us!���`�]M0uF��u�6~������d�����,�>����
Y�fp�1���Z'8�w8^k�!ڐ�?��bS^��W�Y�U����fb��>g�������X7'⠐���h*����@�����c��k(�]C�8^9.Ǚ��S,�گpÕ�����e�0�J*���uue�^��\ q�q�E�(�4[S,���2R��fY�������w�|��x����)«Ja�@����(���3/t�c�e�%�2��
f�$7��3�{a�$��@,�$JnS#�
����$�.n���v�����+��'i8q�4%[ދW�K���{[�K��!Zfk/c�L���<'� ݜ����ױ7�"�D2�V�Ⱦt/̗1�r��W��S&�p�|}'�9�&��(��Uڥ�/;O,��B�`]FN��Օ̤'.y+ԀZu(��b���Q�O�&L�G�ר6�Nٔ^ 9��*�c ��wL^�X\s��Yj eI\�~��3^@��[���C~a,Y J�{�Y�l��	����1�n��Wr��֣FA5V#�
[]��~�"��7�d��e�f&S�%��t6��g��d!����:n��z#�ǂ(z2�ug���n���_|�j~�0��﮳dA����a]/T�n�z�n ��@7��rpc��%���D�i�����I��Y~���s�u���?��:/���)Nb�#1�+
5\*���2(!�+�@\��Z���3^�[�n�<[��8W�W�eeYa�SK�C�'��c�e���ʬb�+ͮ ����;��;s5���D���+sRVb��q#�Vu�#K����X[�������+U稬4ðp�� ,�Q��!_��}c�ǣ8'^ӯ�ب5�'�R<m��Y�$��d��M�"�l�=)���ܸ�-Ob銍o�g��ԛR6�<��f�Ư���'D��,V��<aX(^��c�5��(U���i5�\�W$�q�"�j�̀y�)�j��s�8k\ѽM�t�J+�a�J�kR�d�l%���:��Ê61
����B��cFC#e�Őn}��
%�X�"�r��qr���e�rL�s���yS��< ��ڍ��� �
w</���.��*_�{|:.��(K�z���x[�v��9�D���]N��K_�Թ�Etk[Ǘ,�*'z<���v�I$K������Жi�Bf�&订k�aF]��T7�����Z���XYaf\��ŕ�?ʊ�,l�d'd,��^�K�p{s�o��]���kg��\W�<t[���n��߹�%�.�E�_tD�1��]B�v�6�`9�°������%/�}ӐK�b�xs��ϣvs'<6��%�e�W�Εhn���D�>F��h��(�]�Gm�x�8��N
c��-�ԋ��I5��B/d�i�2�ϊg��lZn���آ�ڑ 6@ɿ���nQ�}tLX��kT�ݡ�;R_�w��!dU�UR�\������b4��b3c�ʭ���H�8Ş9����^�+)ݟ���sF�9M�=m����ȻU�S�FsX�4��<+�I��f���zE����P΅4*T���!s=�kD�c�c��a�WIڃ��"���:�G����W&��w����po��C:��8��#刞�R�5�(c�66��z�E_�<��V�o��:�n��\k�5w�(��������rvr����z:���h2��;��������++]�S�!r	�!�y�}־���Ƃ� -���^�E/���ԕQF\��2ˌ�M�����o�l6e��LAɅ7������*��'�=��d<�Q�R��K��ƅ�zf�?|l�,���9~	��6/d��e�z��r��u��]��]龴!��\��>�5MJ~�/�OP$U���_�z�h�졉��{�+���;Wc&t.0S|�,���<��UY�͇�X�ls���%&Fbo�>�I?^�K�*u��W��,+��+�|rE_�AFT���>jk��e⒢1.r�`�;)i��|(��\�`-Ӄ��7Z,.� B�p�ul���u%����m�rIФ`�[]���n�I�j�sS�L �����R�ݍH���Ui�:i��Lr�P�k�
5q	Me�	^?pno�l�R�<��
{q4.h"3&#�SU�|2��T����t�b�bl@C��Ҹ*�˹>�k�"�	�q�1�>�Y�͎��a �F���a�{h<��r6�J6�,n�s>�"�T�ry>���>�H����(^�ʚv�J��?>���}�V�}Q�Vdp�S���j��ޖ�~�5鬭Jg�+M(��ť<{�LءmooO���o�o*`���g������.��S�l)CIS�p����ρ�[�\��$1�@CHq.Ӯa�4�M�C�E�2XaQ��ReUTF��ğ�zU}����1l�>b{Al�a���5�!6��(�e�`����]#��Ì@��_RR��0��=e�!��3$�����,�m��J�$�=�Zޛ�c��]-'�ڔo�h��M�g=*�N�Q|_�a|�4�+W�Sge�=����<y��푒�R]rT��O��^�r�.]�>G�+{d�C)�r�ݮ�f��}X�P�D9}�5��q�.�ހ�f�mL�[V�A�q�;�m�[��C�Ey����1B�V�J1Wi����塙���"N�X"�Qm�YSs��]��Z�/�bU�+��5��S���Z|]�Y�RI��E�i��1ύ�jV�`�eY�ɕ=I�J�4�.A|���L�<y�ٹދ��e�ρ	��U�D:5(/U���7�e1J<K���1�I�1>�p���S( j(��nG6��2���ڐ�|('�c��3	[���ޖJ�*�ͮD���yrt!?�g����u��u�AQ������&7Y�2�nC�6�rc�u����G?��%2��ǲ��%-�����|�w������]�X�x�+7o��Ζ���we}sC~�����h��ƍ����k��|R�����rqv��ւ��0�<*vXE�����]����>O�7z�ϼ��p(ۅ%�5�MI���e��p���{O=z����+:�|����'G���ɀ.��}����n`1%�"��e��}��5g�\�\d��W1C�sn
%ue+��Al<��+x�b����S��ʲ�P�z]�T�8�h��=�kZVm�[M���OSC?�(%݋c�6_�(p/�2w��&����Џ^�M� �<�9����%?��K��~������״M�[&��[�����1�AAPi,X�q�J]��k�IK>VK�+�.9��f~43��@�G�U�k��Z<iJ���R�]{�k�+YS��&��V��k��I9(��X��K�Ӱ�[O��h�71pq��&]eο���:�03�@�F�Vr �L����OS���t↢�$g�K,���j"�Q�G�d;���8��l��υ�)T�\��2�>a�M�Fk��l��ʍ[��]]U�R�����HNN�8Z�r��]Y__WaO�,�{��ɧ���;T��6�9���C �Ln�mʫ7o@	tegsUv���?x(�d*�'�1kZW啭���TTx��O����\M<(�j(��t�]y�ko�����#q}�S��ݐ�FC���Kmm]�I<��^�B��vd��ʫ����#9�����@�Gc	+x&5y坷䷾�u�?�.���P.��Z������o���ȏ~�C�7k���:<;����w_��7o��X��_�{>�i{{[��[����� ȸ�̌���Jx�^�b����ʕk��;0��!AYӽ��QF�l�U� ��W�U/�Q�VB����d	���#"S�A!���bIx�nC&����ZNgSib����Ǡ4颌#,�y�ID"Y%�LD�k��v9��g�b�O����#�����[/d�p��
Q�m/�������h�(�g@�vK��ܻU3H�6��GUmc>j|Z�fd3u$��>�T��Z�1�j�(ߨx��F蒈�f���KV��9�
�ʧ�A�P�k�QJH$�mA`��x>�Z�S�&�4p=��C<�fő��'�hUהI���U�Y2�4�@p�V�liFe��@��=H�6}s1��i�<����R�u:���"մ)aZ�hB��r�F��s�|,��D:�c2���볜N碝԰Vhpq\�&�%��Mm��Y�	t,� Q}�ޒ*��I��E�P珮?�o���L�g��T��:PW�a<��9L �O%�̤���؀�!���dxN>�Z=���u�b���8#���ٱ$��ͪ켱+�- �j�����#y��C(�T��7��s�J*�].������1�斴�nb=�ݹ*�ɬ"�Y_��ϭ&�������y˵~tBeUdcuM��J[v��%��jw�һ<���mElT"�[��|9w��T��)�~�1涭)���~�;��g�@1_�͝U���w׶��ekkM��[�J�����H��-�dc�om��;�#G����ҩ q��۩�&��^k�?���D���oo��,�Az)��0�щ�w��-yp�X�FK��r��V1�:����.o}�m���������w�����R�ua�U�������zC��[8��?�H��;_�^�����敼�֛���O4G�ϻ�ym(��t���K@��9͆ƚ27|���ޓJ%�:�0�d�iBS?�x��{0�Υ�;UD��k)Rj�Tˑ` |��'��.P�[7a��c�M���%8^z�;K�`K�r�EG�-+�(uG+I8ݝP��Q�LUT[3Y�*�뫒M�R��f��t�=Y�.7X��H
�N��.n��,E�yV� ��0
Si��9ΗͪP��
�80�fK��k��B|�V>Y��肷v	%�V^����1.Ԝ�=U%[�E�q B�D��"W/$K$�P� �1�5�RoU�K�P=���c�����X.�	���!�.��ͪ�k��&6UKb�����H�a$)K?�[0R:��:�;!X+�+B��h��1M�n�:��J]ƃ�a�,0cV��ҁ�H�<2���B�H>9�Z߁$m��f�٪v��p.= ��nu�$mo�8e�$�,�Hr�X��4e��M���P63\�,p�_E��*[�P^����[Zbrѻ�G�I��[���l��r�z������'��ߗg���<�a�ŲVS�	 Ԛ���r�����U�m~H���>��!��L6��e�܄����%>�및9�lv���
ƌ�7ץ]��@�Ai���hu�Zͤ�cc��je��ݐ��X���ěIp�խ}�M O�emwCN����ߖE�"qcK�n�.��9��|(�d$++X�"�P�w�
���!��9_x�j��ػ���>��T����kkk:w����{������Qqp�����������U= j܅��Z��j�ޕ7ߺ#���i v4����c��`P~�[�ʏ��oe1�ɷ�y[>��3<m]q�	O�"d�x4��ߖ�c�g�[]���ۙl�r����7�����ō��zT E��`P�
c��Y�!滽�%��@�c|��"�^k��9��7��{���٣�X����[�M��s>{�	cUE��sW�L4]8�ꁉ'����ŵF��|�����%}xO.��O��e2�{UWV�s�뀙�4��z���*|M�Ê��K�x�8��yA�p3RmU����$�q��-�"0lC� �d�9,�6 � V�l�Q��r��Jl�[�E�¹����t�� �z̏�5d�` cn@(A�|��QP�s(�:�L{�N}:W4�g��"����	��Z�s�x>�IއbɈ�p� (8s�ĖM{��Υ���!cq:-w��'�T�P��7^������ �EK%J���{��&PÖ�#��g�'�)�ܿ�˿�ӃCEZ��+�0�3�8_5�5՝պ�zcKQ��!�8/����SY�9��
;��-&��.!�b%7a ���b�..��:�a_��h��Դ�9Kc=T�w
�;�B���5Ĳ?��-�g��&=(����Aw�J�2�Iʇ�E�K�����lDMYi��~���K3�jE�.���B�uT���?��:==�d,��/��p�ލ��G�U�u�Hk@�T O�>���c�܀ �����.���JK��|�>�evٗ�?�-\s�kocC^{�-<���9�Bm�%�p�u(��;��i��&��(�%�nSVW��ހ2l�`���޺4�~j�t�:�������\֥wܗ��d&sr C1�5�{�O`X<����<W�x�Y�3�����������gR��8�`�I�e�H���鹬�n�����\�&5��g�ƾ~���)Ce�X��+� 	�C��A�z2<'����"g�?����ɡz�TJ0�Ր;�+2:I1�U��4v�:�`�>�N{Ͻ�{�л� E2��R�=Zuv���ƿ��)���d O�N0O5I k.��G��$i�hE�=8���2�=N�C?�3��^���@��o�N�f�/���\Qӣ���qn5�Lx�'��YFy:dK����F����h��ƹ��C���O?�8W�:� |����h5��S(elxn&s�������p$Y�[`sf������;�L���P��V����c�P��~���W�:[����k����f-��U9>���?���*x-!����bk��,P>�] �j�.g&��{�KI@N�UY�AحWd�1Oe֛A�@�,�ڱaa)7��@�M��`E��h���b ݍ-�U(ts%��g��c�R1C�o�R��Wd�]P���>�r\��{7��m�=/cmDg�;�)��Y
����s���H�WW�h躚,Z�܊�Z�����Ŵ֔[T�D�krĊȓ3ل���F����E �����r9oVp��o���	xzHk�k��S�BH�Ԡ|���B>��6P[��ᲳӒ`h�Ay�8����-`�L%l�%#¨c|�Sh���!�N L+��ii�ɍ��,F�>ƅg<I���
х��Ɔ
���ܹ�8g����p�`�y�V��{��m�|���Ԕ1@��H��vp�cy������L�ѥ��n���5e�w�������b:��xfa��zck�"7�x�<�A���֪zM�<���"�>�1�ޒ��59��謯Ȥے6�٭����L.SY�yC�#(��u�+��ڛ� �9~xO�b}���𳻳�h��7ߖ|>S��^��Po
��nhЍ��򳟽���K]��Vi3+�y��w��,�����)��#Y�XuT�������l�ۙ����f	3�	d�%r���IVcJ���7�02����j|����P���T�������zahh�1��<�KI�'��c������[�,u3ɯ�4<�9�֯>} �ېjsKr����O~�Xz0g�D>��u�7��p�1��O�S��D�7��/`,�X�ST�j��֪�"���p�J#��Z�֔���(j�NR�\�5���4�{g�Z�::Q�r�:?=S ӆ�j(asQS/3�Y��^
��R��o:�V�Re�	_�@t�%A��WZiF��âۀ0Y�><?���E�߭�u��Dbx�b�r���M�Mcـ�&��h$�؄0�������&�¢d��Io��!�@2�߆q�
c!�d8�b�a]�.$�P�|ݶ&��P���*��X�9,���ܖI��F� �4,�z��݁5�TA�Z5��M�]�N]��ΪT;���<Pi���ͪBߥ!�%��G3Ғ+ k���"H�q�!�k��ly�������P��:�.=,�6�B�~�_�|��^o!&Y߂��� Ɠ|A�ޖ�EO�Q*7wEj+��d}
���{]��TN�j�\��\ج��� 93���ږx�
$�E{QJ�I�CF,�@��o�Bs���y����;�Z8ce�#M_���8R�9�;�pi�x��P���������=��t>k��Y������DP"��ޗ��'���#nE��<S�J��ve�����`f8�%��&ƶ��V����?�u��ܺ�+��H���w����g�1�ɚV����ɓ��|%����zK9��Νפ���
�K,��5}�s����MyL&�$S/��Hnk��M�ݤ��P4X��Uh`�4sJE��f�ψ���������<|��T��D���/aTb5`tU��N�d{�	_�0n�E`�W�҆��}�P�g�%��3:m���~QE�{�`��p�Q=�_H�]W��Z�d��K�[�!����S���s���]��wHC�(����y�&�s����t���lMV�xև�����^�!�;�Ĺ2��4�l����*-S�L���ǵj��oB������ʞf�Jr�3ǁ沌��J����jx�����B\���CH�Nz������l�u(Cck��Kp��7,�������� �2i�X��tN֌���*-qwY~\�L�� �u H,z�A)oX&3�2��չ@�K��y����9c�ЁL�Z���FA�
avA��f ���e�4��dП�CX��t���p[(^(9l��E*u ���H�t2� �}�
���iA!�'�LH'���(2%C�݉��}&
!rh�~ʙ̜�㿕��HJ���RĂ��qt�c�b�q,Ӳ��Tp�@�㹎���X@ ���P$@�HX?��w܏��:d>����-X�PT۫2�(�JGn|â�{kJ�5¹I�P�㹲����[oHB6� 
'9j*)!*r
������f ��P; ���o��o�a{);[��n��>��B>n0a�p{_�?����]ZV<�"8�����Ɍ]&�yf *��}�{�t���}�{��dx��0�N�5V����)��{����/��â��6W��M74?��㞬T1ߣKa�\�5�X���!w�"'�����̬��P�H�r����d�N`@�e�-���zN��9��,#�������D��ʮ"9���ϱ����U-O`$l`�I��D��M#1REJ���mP���I�(�:��rCq�2!�b���?�(}C�3Ě��nlɎ ��h �x�	�k����_a\�!|vp�F�Hbȉ@��1F�����g�{]���ʖl��M�c�r�W� �jveߋeFpL�.���3�Y�1Y@<� ��{�AMv�D�_�Y�j~�q��)J�44ʭ�܇���}�|i��$+o�����s���\f��*��n��\�����5�\-d��J�����lXP�k+�Z� ��3A\���:^z�+�g�?�y��KZ7f�	�a�q�hm_��(7c�sY�B{v ������
!톰��*t[S7�|����Kd�ڕwn�",�&%$Pha#�2�do{hd��K���8��ضMI[mI*X�L��Q�Nu�E�(�n��B2�'�$�]iפ���a�kV��f)PA=m5��}�p!BB�jE-�6�C^�f�M�M�ƍ�4����@1���#1n2*
�6��[�K��gf]C����������&���wߕ��Rvoߒg���3���M�r�k��������?PT: ��"������;��������d<��
s�C��Wߖ�7��pp&YE��Is5���\�7�[���\B><8�$�g�Ϊt�UX�k��~K>��ϵ+�{��I��綻-k�+ʒ4�b۹eq�����ּV��70?�{hU����L爙�DNEK�藊���S�����v������V��g{kC�0����^`-��`��ｭuY��o3VʵFW���<�\�u�����|���H9;�"	5ƹҭ�Y�fBW�+0����ˤןj�z��[Ե�zyvr�Huփ�r2T45��*My�옅EZ.������C�U��RV?{�\��-U�DUMlS�/O�@�@�������X�-(�:���*jͲ�{��ӭڀ�I*D](�F<�j����Z��'�9%�3e� �U�ʝH	�'�UP�4PÐ1�v��[�`6� �B5�2w(�V�l������o�u�'Joɺ�f[������4�9�3<K�=sl�X_���Z�h�s�!bo�H�m������a��0驳���\W�)�Sm�s-*;|�oH#��O��;w�ʽ{+/�6��������'����FC� ��M{&Z0��}�����Mc��ܸ�+��Q��=�R�_�#
`OV_9e���"Z��B�wdM.�	Sl>O�@Tj���&�0F�:���� ��c\���B�o�hk.(��M��w�#�~�C��H��We�6؝W^�w�{C����0�6z�&�`��@[[r��-��Bx5!Їf��A�om�J}o_�3%3ov*rq�1��!$����n�)?�H�%�VU�!g�)��My}[��/�AW��p�%N�
P�;_[��?�g��?�;�^���2v��o�`��䬥�d��0k-���P��z�?|�l_ܠ�d�;����ʿ�˝7^����0>\&5^{SnC93;��[�� ���-9<<�ݝ������k���]鞜�i0W�Ԁ�g����VC�@)��O$M��Z�C9c2���qkϟ�>���4�0�y=���R���7���!��z4�H���r�?7F�u��t[�ߨC�Fu-5��Ø�^nT׃ջ�}�.疆!����c�q(���L���&��\(�F.�ǚ#��@�{2�غ���40<���Oe����d����8c��Y���#B# ���@�#(�Z�lF2�aoLd8��y�UU�I~�)n�F	��\�Df:�F�&3��������C<R�C1%Zu<�����Kc���.��rc�2�S����m���2�Y�DŖ`��<$:���]@Q�jʨ�kW�t�V���z�j�ٸ�Ge9R�<!ဟ�<����	MƑM�d^��G�y�:X�L��+}�O�ҹX;)6�|v�%�ؑ�1�%aq�uݰ�zU(RX$=�V2�4�!,>���zc]va�_<}�׶�I��ŚY&1�w �5�'DK&<#���H̽�=����sݨ���d�b~�kf���Ho3���yN�?=_��{#sa#��N|�%;^zŋEik���PQǳ'O����*����Z��
5��S[Uݬ,S�c7L�.�W_�����S�����I�v����i��2��¬��oܑ_��WRR�{�,Bl����[�z���g=Hy�&���L�ro����]y�$�y ˲��)��@�~���z���i�oɃɑ
M&�L�UiuW������_�� TI.`�_V�FcGFY_����+���&>��yS~���R��ق�]o�q��E�p��r|p��Ϟ��J�ڎU��jj�|�%S)s�}�䱴:]�����G���s�9�~r.'@J}(�*�׾���q|��l�Ve~r�4wd
`H��> Od�ƾ��D!O�����Ƽr�������˺�\Ά`@�] �l�m��ۻ7��O�{J}�l�ߑ�����8�t�P�3"$&iA�������_A�~�@rs9}p�(�J���s�^�Ž�r�]e|&H�ۍB�{�cj<�M��r"�/
8�S�������އR��.�x���ǵI�G(�J� �=z�5��7���y�al+8���C9�5�^�)��:�^
�g?����74�L��FѢB���XEe��1����T���J���r$�������j��L���sf���{��t�4�k��\Q�/DlK�/����xW)Q�J���s���@�^���J�Ť�5�c�=#��V�l���9Rv1&#a*��f���%��j��=�:0��Hgg��'������n�p%�'Y���R�; vf�gs��ikX#y�1�K����ZK�޺bɟ�}[w���`�K��@f�+ՂB�y"�k���,w#ҷ�M�/��ö���F�rd1�"?���h�Q��q���~�����/��	Ppvv�I]��� �����"c8��/���B�D�j(
��ĭXf�h���K���џ�Q��l�eogW����]�b�Mc�a�^������|����������2NeлT7�ڝ۲v�L.�Z�q|~f4~l7e~��-�������w���{�1jui����5�'G�3�C��i3��IM��;����b���-�<=���-!oBq��ٖ��@D�ByJ�����k���=���/��g��H�Bn�vG�=Q��S��րth�6���QF�q�3��?*�Џ�cU(���U��?�wr��=�Dۦ����c�Z^u��|���*퓟�/C�у���Cy��M�k��:yj��X�6����)�L�ڐ�)�`s����zR�\��U�اm�H�&y����顬���$���@v�z�\>��	h,G@ߏ�G�H9�%�(��b��z�G�ޗ5&��n��J��9�γYX$X�su�>�j��qYnD��9W4����B��,+ʡP����P��1�%�֞��]*���d���.����M%���'+�o棾D��*8Ǧ
��*�v"U�I��>�V��v��[��47Eɚr�<����Z�%A�$4��lc�;��\Ÿn5��tm�j(%�j�Z���$�g��)y�Xx�/�Qc�c2v�x��iH�]5S ����0R�/Lr�ђ��Z����Y�hs��dR��5�U��x��9����6�ky����J���KM=B'��I�#]'�M��6����ElMYBSp\W�!0:S�9��AC0���#�$7"1�;�Y��T*sk%�� �?�k��U�H����"!�{l��z�d(,�\��3�9cwE��"UCT������X8��=��O��p�_^@�u�Q�`ٴ^D]5�:kaܲD��@E�2>�H¢�X��?���G@�M%� �+���؏>��Jvܓ��u��������'�~,��z?��ξ�6�dr"����?�XN���5I��2崆���3�ֺXOT	29h�v��g�Pw6ߐ�������@�.�����w�&g��������'?��|��ϕo����}S���'�7oȓ�Gr�;��h��K��ew�����Mа�O�W��܇~����⯿/w���ƜB0��3l��k�)�<���d@L�PbU��\�Tٺ�B�B8Aa����c�B��si���e���H|v$k�P�˱4�@7���s�*�iĨ�T���S�f���w��=9�/�` �h,�2�=�=�w|�P�� ���l@�N3Y��68<���X�XG4����"��nG|;:M0�����O��3��4�� Ѩ{n:SNb�;��RcV�0g�B��b��r�g�qɀ��ĺ��f$kɭ_,y��c��<Uv1b>D١�v����5+%�k�Wg�!C1�M3$G�� �0���B��"B���Y�
��@P�Oa %in?IV��#�[�=l��G�V������r^�I���*�;֗rh�SP,{`o,F4,0�ܲ���5;� ����,�H�%��^[��s]�m1�zғ���Jx�sB�0���8jm�b1Ř�bͳUo�$�=R�f�\ۊ���{�Ơs�f��k�{�%�|X�p܉����Q��5�6�B?Of��C�
��>�1C��GJ�A�ͳ�s�9"}��En����L5�Li�6�ZUI��Q�@��Թ#2C���7w��/����3�A9��e'�V��m�<	�A�Q�Mj����F�[�r�衢�H�bby����_��\������=,�XKd��$*����L���H(�\Lz��)����P���' H�2���dP�IGkp)��:�&o4����"$!H�mpY�K0�g��%l����"C�={z$�ˑL�U<,�����_Ih��s2�"��`Nf�ҕ��b��f����OY��1Q�0�����'|���?��m����ӏ�:��0�Y�=��(�>�9P��{�ͥ��U����}I؁����_h&tDD9@i`�O��f@�@����Dl��z)O1AB�y(�32o" 6�{���Ls<�h*0ZokG�$�4����@bf��t&�l5�ڐ^���\���9��@�꠪n�(t|��Z���������P�2�Qqг@�>\�7�7_��-�[f�7�AX5��Y蚼��x5��d�����c&p1�
�wj��a�	熜��\ϳɬp#��L����4,�{�統�-���Қ,��R�Ҡ�[]ښf8�5�1�Ps0�f�K%$�.2׈=-ܕD�i2Q@6hN%ݱA5��s*��eI��ͬ�n�i��BaY��;��JT�IQU][�X昻1�0��4��H\�/W~�U	Cz�&�+��J>#f���>�?k�3O������)M�hj�%���w����0���!)`� <����2�SvA���S�:c�{�믻�(��NՀPT-�=��Ϫ��f��5ø��KkHv���al7��TK)�eq_�i^�T	c*U� [0�B������#�d�W���~�A��&r%ӭD���ZD�Kd��Z��U�v�Qw`k}JWRE\h�)�3[�1�����S]@�@�<}~�M����ƶZ��'G�rtz$ǽ�f�VH9��[�x�{
���:�8�_��X�f��>�ാ����Ca���@IR�F�#l�秧2�f"9������#i�Y��j���Ǉ����c�7���!�Cl��ؗ��9����O>պa�U=���E�jR�̺�0q���|�>х�V�t%s#��c�ި?�����T�L0���[#�	�	J�	� Z(�O#<�f��ҟEl0�� {���?�VJ#���D*���]����Y�e"[�`U�ZWŚA�N8f���N�Y`�����^�_P�J �� )��ؙ�1��jW#��H�m ���U)8�n9ESr'�|H���Y�Dk�w��%�Z;�8��ZK&���l���<��:������dx|	(M)�ϸbܩK{}Ud<�d:Ѧ�i7%ߵ=s��1��ず����uq�ͭ�]<��wI�/�(Bȯt�@�-9>�bS�`��@G	Z���������CE3�T�����6�ʧX}�*P�׻�>�o~��՘H�6*<���03�xN:W��\K�d�Z��Z/�ؚ��8��%՝cG-7b��f�-ڃ�ߋ��fnr�^�T�NMD�4�S\��_6��������J�ʮTZ�#\s1���p�4���NǓb���e6�����V}�\nIyl"B$��9��ia䭮�h=��A�\�e^�Rq.�X�bI�ψH��k��ܺuK�~�ӟ����*�rt��|��/���+^zq��^M5dd}o�@tq`�ҭǸ�'���\�3"&���j�h�;�x-�H��L.ԅ��C�V%�1��9������>��%��M[��`�P*1���)��+,IB[DRoQ@�]��?ɠ�޲mu��"n� PgP4�X^�����%�ό��M�#5��Bـ`x&�LF�������FL~ �n�65�c��zg�r(- ����
/���+�~�ڳغ75+m��mb%��tF�	�$�̵��{D��1��LA=g�:�5��I�ܸ�)$C�}�)P�۵��S!�l@�]�=�O�Φ
�PƘ�	�C��pC�TP�(��!4I+��xx�<7˲rJ,����R��-^MF1�;��c=�FJK#�.����+\}����5(��!/�^je����?��wv��Z�Z$X�Z��D�Ԙf$��7��Cy��1�m�/|A��8"Y�ݑ���2e�X9?L*LE�&�؄J��we��g�;�)鲖�zC��M�S�r{�L㝪�*U�.�w9����>��%B���Z3��*�T�:*ۑ�5z``�(�F�!�ͺ�)]�>������}OϏ�E%�f5I+��Wi�(8������bͭ�־p�]�B��0W�*bݓ���4���C#y���Xg��Q�GD�|6V�L!TS�~����q�al/�PɭoV��bZ�Ey�IFZ���%OU�j1D��4U��X�Ɛ%(��{7=�c��Jv2�*��3`Y���h��^����**���*��iwdkg[���l�*_���<�lp�<���K~��7�(��FJ���?�X�h�[g^&.1�B&�c���"�ᅒ�@\��X{�F�B<S:�jLE�J���imt4�[�031��B���h��h���1�g�.*1�Dp�]��\�p!�?�rj�m��(��\���}f���а�7[[@އ�̘TJ�1jZ�ӑƯ�P���cĦZi�F��i-]^ix���퓮�aY�p��@�$���ӕ,9C����7q��J��{�!EJ�Hi\�����!9�6���ڴ=H�[Hg��=Mm�0a6w�F�J�Ad�n{��z�T"�s���t����fS6�KB���B��R:նt�����K�ʤ�,�8$�V����^O�e���샨F�(�֪4�k2�8��G5)�G����s�h/�g???��1���կ�s��w�nH4;���{ku�	O�Q�h0�R\C��򶦧s3�JgjO�;�,�:�I��+�"�`�\�<��ɩ*��u��ݓ(�/// ���ﺎM�m���;�����HP�F�Ŧ.�D���e^Pz�~O��~U�9C�h�]Ơ+U-
\�-��"V���.X(5��N�y=�ᥬTa�y��O���T�;����Pb��:ka�\�Ü�`Y�ݱ����3^W��lFJY�ĸ��)�VC��1��k.�����D#�-����vG�4	<3��5�f�l�� �TSR/�K��}�7e.�[?f��1�j�+ʦ��U�65�5��#�,�1� �ʌ�k��s&�e׭��m����InMU�]�\l����vңg�H*T�:#���/��%C�.L�W\����Bf��nn1���g҅R���+0VTg��a���
"1��Jf����f�+�� �f�X)9�a�'�h�nK��e�ز99>��G������ɒ�|�q�̘t%�T�A�!�:��`�Senq2u�J�/��h�@�L�A����P�&6J��"���s]]���5���%��Jg�HZ��-Vu��l7�g���0Q�?�������eHQ�m"UC �7�~��MΥY�4����\V`$������G��&��F��	!,3�U��2 ���T��ZQa��,�݁�k�I
���Uk�T}�U�z�-5�/��?7���L�I績�<�d�Zzfmϸ�6֤���̒�(tFx>$9 �/��֒��c;D�w���c�K����.��,?N1�pm��Τ����:�0�ų�:!�җ��C�v���P���?��f�g秎���eq�cK�#D/���h�b������p.��a� �Ř�fjSs3������V�y'�]�(dG��ٹ�'�_�zFk�H��i�0�O��J��������I*��ԍ�N̝��#4�0��dy?3�Ӱ�	��q sY|?�<5�N����+u.۰V׸�s3��C�N��?t�Zl�a���Z,c�{����"֒����Ȓ4P�(��	��z"]ЬN��ݘIy!�Ɩf�O���9��k�%E�Ōa6h�(Gs��ҙR,#��y�+��lp@z� @�	�����3��Y�f�F��X����J�4�Nȇݴ�pq�李����/>���ݸ��V������0\�2�pï��L,13>u~4��{�����R������!�u�H�tB"n�V�����%K��SY��������b�����7�яΦ�澣;U;�P�du{G��ZU��Y2�0γ�ؔ����%�W׍���X=�X�Z��w� Xx�H7z��
*R�*���4���H�$H�%/&v+r�����{@�Eu)s��ihy���M��(��ؘK�C�Lf�Ғ�^���<�ݻ���G?���j2�;!�:�jR2 �y_拱6H��rS��@�A\�K��S���%�%3c�.U*4�dw��	����t�0\xϤ�d�PBWq�~��`�߄����RI0?�!WR��f]�"ʹ�$�W��b��c�s��_i4O�MI��j9χ����?;;Q�&ۡ��]��T�FÉ*�I2���3���mx�7�pƠava�g�Y������V�JM�u�ɤCb��ۀ�?}�8��sCET�l�׈7���3���B�㙪@�٭wq!+{V��d66&	1�r$�(�W��fW�κ��T�k�s5p�+����q%�D��Wf7G��PZC��֪�lt�g�N?LS�
��h�������i����+�%�a_.�J�:g�fm��'.t��(�/�� �̬3��EbD��S�w�W0W\��֋���3����zZf1��-خ��!�L;AեC��{uN����r
�co��iA����E��MR����pl��ĵF���O`Б]rϤQ�����7r��>)_4��4�[���@�q��a�p�Sf]C܌ss�{�[�iL�|�����3����0�Fj!'��י�r|p&��>�P���P��L	�2L�l7��0��`<�\�e?��re��p��/w����~���֛J���z�Uc��i#�L��X��+��&�r$.x�c�u��s$n`&cN�4�lJ&fY�fU����B�,IM�*b!�ӄ`
4�U�@D�%O&c���g��X���vX?Jwz��=�+r'B`�<��$Bo�[�;9R�;�:�0���Ko�IH�%�0�Ɨdi�sA����Z��7��//�䈙�l���LIV���ԝMW�j3v�՘��!r��d8�M�P���P���;Ӓ�`��1k��M��@�{a K��"$Ȁ�����N�^HּIP��\�!d����eY��'OKĄ�d�udB�c��hГ>*�^^�<r�.��ԘWP'�݃�?Υ� ��$��]�����K(�<+�e�J#\���ω�f,r�+u1����*	�p�]�`�kx:`��T��x�P�Tݔ�C���h�9o�-	-��-V`6�����u����b=1Q8�4x�7GPtշP�XS>OR�:��~gKN��wZ2����+��6� �M���(������4E�$I`��pك��P�g̾'b���=�U�$� cS�^���S�[V��t�>�H�e��̀�5]2�~=�nA�`,�L
�51_0"����(ǤaL[Xo���D�/�`x�3�_f��
ńL����+1̫F�f�Z&���<jT�x#E�D�FbF�d4������ޛ��vVU�su{�ݞ�ܾ%�$� !1$>���Z* <�����+_a��S�*;�$6� ��ZRjB�(���雛��{���ս9���������{W~�wr��gﵾ��َ9�PS�����.����n�h��p�8J�����^'��eY��U�(�U�Љ�`���9�}�l�9�6����tՙi����Ō�+��|�(����	�L�$�unC�G�F\4��{�;�eC�D��Y`5@F�]�����a!8Ҭe�N����SuH��@"�}�1#�U��>���mC�#�pQ&��}x���lmhv�JX�B�A��>ϔ�	��Ad8,˟MI��)������,/���wc%V�Gɂǁd�3 �3���D�@�nl�#G3F��񹚊���	��y���,Ԙ�DU�R׀������eM�{�?m߈�]��#�aە��Y�l+���	�V�1�<�����S��U�>��O�%�@���3=�m=�p���C �{�q�H��(�55��?(EB�P��e�xCuTb�ߣD�~'Z !SF_��q`Y=��P�7,���;�-]����aD�wa����l$�
�O�e���Ն;4��2}��2@x@~�y������F8jB ��(����q$�fk�"!�]�`�Y҄�C��f� �2�Ab-�K3�/n�V�9+�"��ޣ�?�$5R� �ip���K'��]���s����Q[����
�+��X�<��R���O��R���螝��.� �[O 0
����(�_���ϺO�.<� �Nc�����4��f�J�e�u�4 ibf�Q-���`"uO��6�pA��"�~#������rWW��v�3�q&�!#���k��{��;��h]� ���a�
N�Ơ+���P����7�K���r���:�]"�)����=c�Oy< �}�Qs�q�6`;2D%_���x��+�U�����švC�N����:˾L��������Tcf�|�h ����̈s�ۀY�jEc}X(v�@���eB���X���:����v����8L�C��X�F���>�	����Ô)i6��PgIm�F�����,q�`���X�cd7-����:Y&�Z�>%J��b�c
�Xɟ�P����D�K��_e����Z�y��ٻ�d��ӯSu<c?�N�c�E���|i@��؅��.��L�Tע7K�}.�77��s3�0
�G����>��D/}�N�*T�$���2eI�5�=D�0tmݱM1��L!�3�_
}*zYɘ�rJ3�����֜�$���p\�A k��LD�j�n�h�u�3�����&�=ʒD�D��ḠL`p�c="���I�Y����\��A��[�l��f��@O�f5T������yX7}]M\����e#Jぺ�85����s/�H�-�����C��1b_�g�l8�r��Я4-m�Vw��˫GMj&|n}�pa��W�SW�c$ñ�	u� '�^3z��'��nu��]Gi�ˮ�'������5���R�K��N6k�{�e����t�<�&׸G��R,J��O7w�������S����24��>���g�����}�XekC-H��h�g�ғ�&����lo�L7��a�=�\�M��������ߝ����ox�|��;�=D�K�����r��Q����dʄ#j�NP��+^n���� �($T[kt�])t��o#r�iE�i�z\t�Ɠ�L#`_k�pa��0���xta��	S� �C1�T�E-����})G1�"�Y��wD1�e��$(�~$�����Hd�q����7p�Y��I���c�l����p�.���	;�Bǌ�	v(�!�ѯ�]N����ܪ�1 z�&jR�x��mY]Yԧ����6�txE�\���8�%d\��!+f����Jp���@$[8.��!!������2��P4P!
��	dC���9�Q2D�W?7�i�˦1�5��Q���`�K��B'3���:���2E���Jj0�qZpf-�%?dj�CU��D�	Dm���h�^7J�$�/��,HI��q�1N����ʱ��9.Hb d-���|8g�ͬ��VY0�_�(Z�3S4j���oE�es�z�x(���Qq��P�9�H�������&�	c*�)��@ ���:`d���=�'Gй&<r�ڱ�-}�"�:	���)��)�b�����bG���|f�����`BR�(�}KA���{=�7tM*��EF%	��[&��bs�����)��ӅXC��+����ҪL6��W@ֱ)�zS"u@��.%�2�#�7u�ƚ�������S���Ʋ�Q Z�C��̙'��P���j6e�:�-�6�}�G��t�����V��Ϯ�;zv�c�O`��+�|VX�l�>Wpx�@�=�gF�1��Y*ƃ A��s�2��<�>dl���/��#�7����߆�[�놳�k`�c�}c)#��hT�T�2h#^�C�gly�j���H6��h�9ؓ)Pz��H�����Oy%��!{9��%���|�c#��18a��1�d#��BΕ�	߷d����`��'�$�|.~���rd�E�I���Z����	�Eȿ��2�P����9��Q�fݭ��Q%ȄE���`���S�دB�:À�D8��N�j2��i�__�y�AII�@oa�Ft��>�)2����H�n�?3�b�׭7Yo�0��H��x�=4s��i$���u]G����ցҏ���Gpz-���qMYi ��r""U�:ЌӨ)J�m���	2��"F�J��:�t�,8L�T�0���}N�\8�C ��1��j*�2����A����Kg�Z
X3:h�dmS`��luQ]��ӦE�����h@~.��#��L\���c(�(�a
4[a��\����G�[����
e���T��h�� N0m��4H�8�lp�N���	��(��y��6�ͨ�~�E�	̜v�)������66��B\�,t�	!��b#i��k	+Ѷ4|i���@o�wx<��xۨ5&,�#ۚ���rq�4��؍f14�H<�Ni����bD�ς:^]�]�b�:g���v�Q���C:��k��d���v�;�`��]=_}n������S�{��������	x�50yd��' |��uLI-������齜����9�ϳ�h�v�)aF���d�z�*����RgA����&93���"�V��5�m1� #+f@T��C��>�R�J�ƕ=��4��jp0��EP��3��(���x>`����P��'_���x�������+����>}��;�=��3�@�vw{�\㩍X`�4�G֚jԑ�2�c^0����P< ��Ԋ�9>@��@�>M1O�N3���e�K߉_á���(7Jz \d-�h2��m����c�4�oK���&�c�I��EM��QJW#
���s��6k�1
�����,�|�T�u-����=j���}���WV��xI��</��G&�1�S�}Ǳ�}k���5ՌU�YS�!���PC�	�\V���u�F*]r�tɨK��5N���PW�/6�,��_֤4�:�����)ʧ���``2d@ꠙ�:�z��d�O6j�Ĺ�L�g= %Q�kdTrs�ɤ`���y����r��������H!��Q����܇%�$�D ~0��I��O�Y�:��s�����lyDd�k>�?yCwB'e	��@���`�H�T��D�C |ȹsz�QK׭���(��:cF�N�E�6D"�	��}Y��S�5C􁾯1���_���׌0˚�%�� 3�^j�3�_\�J��"� u4��49�l�q��� ��l �=͠�l�C<���!�S(`�y?���)��ɢ��ި�鳂���]u��.[�r�-i4�$^Z�Ϻ�h�g+�L����P��{���k�lT/Y�2|Ǻ�[�c�]�JTk�玹�>��;���L�K�����)��\�L���ݎ%�\�j��?�甌WLT%SGmk��̕�K�&ImX&H�4�~g{�@K ��*�4�` ���ѣG噗^�	��:�/�q��{��9.H�ۢ�@��̬0F1�
��2�KO>��W;{Z�+����w���t�@PR�� 0��8C���{�_N�8!}}�Iu(c��5n�]���T�į5����0��Pd�b@*�����8�1��X
")�A�未AI 
��m�X����@�l@�[h���9`؟<���>T�(|�A��Lh6�A�#k�aN����)c�z��&Ř׀Ѡ^_i�A绽��1� +�Y}��'����]s���c���qo];�g1���u
�<�b�#����#"���拐55r�h4���K�馹=��jƵ��M�;��5�wj'���ΐ�9�^�\�{�R���2�,��Zf��N#a@��>M�u�!A'A3��BO�����
��F��F
&��t �f,S)I�W3#'\ ٨'��, O���rv7��+	SC�6�	`�c�� �<��C\ãIG3ąV]6�l�dר2�^k���^< ݵ�x�����N=��@+uϪ#����~&] da@k���H3�u͆���OW�S�W��D���6�����:u�}8}>bO�j��}����(5c�v)j�/ȱ�%YNN��_����k�30E�r��!���|/t����:@�R����|���" D,xv�#H�B�;!�<�R���P����F�pp$��X.)����^�a��}�z�#W�9�c���/ `(�U�:� ���٘x��:�FQ�1D.[���ԗ8F8� "0�M�J6
]��w
B�%�X�}����R'�"6��씕=Np ۵=�"�E�)
�r�U�6��3T�8��i�c���M���/~���&�3z���8��H��vQ�B9��e��i�=ٿ��n� �����G�Zm�ƈ⺑u���5~p {�T1����CCT��
�T���}�NM������F���ES4[����,s�Y�}���~�5����^\ާ�̓�O?!Ϲ�2���(���S,�W���P�	M�HG�-kv�#muf��TF{j����Pg���>�y��7�����lsw���������YZ� ��s���dol�(��dGb52㡍
�EYw����&٩�͓��H�fG����$c�aqYAO6�7(���Xy��'Ч��(����e��1)�&zj4K�҇�P�<���<,�Mi�}l,�#NY���cW�׻k��Kj<V��:H�%�KewX�{uL�́t"=��,�ؓ�:bu�Y,�i�4�W���;��E���6�5)d����m	1���J����b�+k����q$+=W����Y�<T'���fn ���͠F�ʇ�N�����֞8�O�:̾���|'�7���Q�n8���:k�?b9tiS"�O��3?� ��� KGNI�k���t�)��c�m��kD��5��Iٞ�j2� C?^֏h֭]_L���5	��Nv F4����4�����5�zU�<��6۲oeQ�uO7OjP��ϕ��4z���]^6���C�Y���}NL�:H8܊�`Ȕ����Xں�.;u��pi���.�� ��G�`�`��T��&Bߘ� !�3��f�A��}��MĲC�M��p�j�+Q�ؘ�GE���vJ�c]�H_�T }���o�CFK �C���( 7 �4�1S��I?j<6Շ��z�JP���R�Y;��U��o�yDp�8���ԁ
A� 0m��+Km�����N?~��"�KK��c���
���&Y�
HE�լ�$���'O��璘������o� Z��_YJEI����k�5#qow���KHzA)����Ϫ��.?ړ�X�k{o$���t�k�u��q E3��;$`mitd��)��e����t�o3i�|�:��ȼ�������p��c�{�z_��E����Lv{�yg4k]s ��$�����`�:CI6���:��A���������@_�+����-�>3f���M-R�J8()��Ǩ?�(�!���k�{pG��-+��A���=qRV�W$Q�9I=5`$��X���s���	�u�~]�"����Xև �f���-=��4��v����^ڑ@�s���B5�˭�&���N��! C����Mu:�f8�/Ͳ�z�w���@�#��T�k����� �K�&�bqH��pϓ�m޳86ed,%�3`�U����C�dK����O67��+����Ξe�엵�Uu�g��OD�֥��j'���ۥ�ò~蘍����'4�Ԡ3 Z
��	��$�~umE�V��g�'����w���d443�PN�Jۃ���:̺�����.
�x�v������5*հEB<AN6�NS3�t��$	��!˥~B<7<�UC��d�\���g@��h�-Jahg��&̽	d�/(��I�f��!i9����2Z�4g�Xǘ{��8��=�w6ͩ�,ld���91 c����w.`�֔qr#��&[S<݌�L�- 
�xn-{�H�J/��d}}{�`�d#�q)خ����8~P"�I$����� �Y�9�\�}�	d�dj���f�́��� �T���#ه�Ȗ��>�����<����l)��ӣ$�]7ղ:K��W]�9QC��.^',嚴��ޞ� }�ءF��z����J�xX}�p�\�_ȶ:�/�=+�.�ɂ(P�AAg�X��·��C����F̯No,�[N9{��Hz&�e���s������õ��!#T 4��i�9��#�b�@���f��[�� G����&mK�I(�Ey	�O@1b<ڠ���qX�#(Y������OȾ���N�  ��,��N�dA�� T������%��#`ゐ����g���M=o(S�!� c��J�=����(ooq�T�kI_��F��A��2�8�:�=$LFj|�CP�W�o%f�tcF.Z��-�ӏ4��A`���h ���YS�U�C���٥��j�w"0���.���k4E�e���	@�v�I����$!0�Q��-C9r���������`�_��!Q��SP���2=���x���֒:����Y���p����y��H��~�H+�d��!���o�뀈�t����Gi@��h���i��+��<�N>�1�ڤ~�$��L-�,�?R��q�"$��K�f�}�x |S3�CΒ�����x\�,Y�e�IbF��<���
AA���G��>�]9>56�1�9 p�G&Y�Q*D��G�g��T*n�t`�;w�P����/!���S�RǷ���a�Y��L|����5�N�9l���z�s�q�a���}-J�n�I_�|�,��8ν'n�/�}�5��_ [1����CqNP��*	K/0mi���:�5B���o��{����?���r\��w{g3�[MYZ^fo�СC����%�ڛ	K(��:�^����}+$K'�~eYbo��]&�6��Ƕ�ɒfCP�����8~�s�@r�_�;xX��9���P�@�i����{\����'0j��L`��#
t��4k�l��D�G@O/H�I!Ф�Ʀ�
�l�?�.zU͆���n����T^��z����@��#vow��U]#� �F�d��S�ME���l�i
 g�������Y����fe��"�\����Ki���e�/z��;�� ��AĐYV��f�k�Ɏ��{C��|�{Ӿ������$>�SJv��=O��D8�xY�ỳo�����F�d�)�m+n���ًj臂���쭁�M�,�'A���RPU�=@�����Cp!����p�c:���`6�Mܧ��%H��`�&)�l! ���?�k��=n�Չ��;��}�O���,�	E"��=�Af*C���0��bJ�=���u��!C5�JM�S�hԁP��"F�|S�!��F�8f���5F��$j���O��u� ?�H��.�� �C�,@x��/y�Ŝ��8ʻ��`���&�CX���IG����G�
Sf�S�O�	��s�kE���s��_5&��G��)�R��8{f��;7�R};עpζ�����ke��2�ަ<�9�6
�s
�-sB��>��S��pD�*Y$�AE�G-$Y�q{G�.���\�&�s7��1�����0���{�����Q�����&��cӠ��i5�ٶ���G��A��NhZ(�iF�h����f�L��=��^.G���'�ﻗ>G.?��ݺ�#�Ӎ�|��t�n?��i�����J�?	M�ԟ�)!Ć�,
�hN���}�2gk39qtU��
5"#̌����dHZ=�U� >V5��f��蹂6�h-�ȍ��xB`j��S��ܲY��ðt]ƛgfmB��EƂ�<��Q"��[]]�5��$}$ud3��0Ggi���ehP�&#�S�led`"[z�`;�L՘����Qg��:�RCN��ZdZ�Bi=%g�i&�IC]#�54&�0%�� hdpAC^/H�=G`��3J>N��-�K@����e)Ef��O|f��X���������0����J�C+���k���&��f��	i
Q�~e6FT�0�!�hj�`�C�I��陸=Us� ��FV��qQI�{ ���9��rt�tj��X�w��F�N�7~k*Z	Qߘ�.�?@!9u��PŪ��p�\���x���p�I�a9��z�(:�b�ecĝ5�[��G#j!Eh��6A~�2t�۔���ɲ��U�nu�^Y�u���5չYY���*(��#w���ԥʷ/�uA�U�U:^�����J� �a��}���d9��V��95��	&:�W`.0ҡ�]�,�
gLR �r���Q����M��dD��]^^%Q�/�⇞��g~J.��w����8�b���ٛ��#D���:��.˨�>��:1�0���G�f�l�ܖ,�5��M�n�ȵ/�O-W8f}�vD�����8$�QK�`�X��$R�5k���Z�ĕ0*E�*%�B
�N߈"�p�fQ�@�ZRH��R JD�ct(�$�VR���2u`�'S3<0�d7r*:����C��l�HR�`���9�99�M�畦��p��J�!zng�P�8>�
�b�@\F��?p,A����=s�� "�f �e��3�bL#M`�eN�I�;�c����=Δ�t	 ��g�;@�RP�`�$48�-��@��r�)�\T��L3�+&z�> �}�V�##��e;2��#�(��e6��Qt�@��rJ�����6�����5��`�S[�B��F�ꄢ�G�j��	9� ����M������2���K��sn ^`�&�K�n����t�}���e����pA
��_��Q�)K�Q��sU���:�Ӟ9*:Rz�� ���)m��!+[���޾��w�ϥ� ��Mޢ*���&�~�C����ܕ�q� ľ�]y���YH��L��`��T8zF,�Sв2���9���r4�����+�� �=ڿ����g�,A��s��>����g��;�9��#�Ϡ�DEq8}��+��������}gk�ߟ;�(�;;t���QN����h L/��A���⥗]E�d��d����:��\�� ������`C��@�q�U��W�	��)4Pp@��Y^��U�0'�cC߻I��O�n`��@C��&KK�p$�a/�!��8k��#�0at�z�q���fU�%�؄�ۚ��(��Q�B��â�F�A&'=g������$�L���f����'��;<�Vr&AJPcy��u��A��\!�g�)`y.��ɹn�MN��AR�2�1����P�)F�S
���=	H��<����K�KŐ�	D���ӡ��=�"�˙)�0B����9{_ߕ$���W΂eV���P�,dB���l�ٔ|�1����Q�>R�^��,;�H�u�Q�Y����7F�l�@���E��~����"X�87e�DJTJ\(6�u�BND5dߠ��4��3�5zb�<�[c�C�A�qJ���م.�-��� =hn�[XY��VIڏ�aϗ���,�)$��Yf������F����i�P&�'n����;Ϯ��;�[f�6>f�cU:�dh�}L�&���H��\������9�۞!��D=�W9^�9���e���Ži�]�[��]aׇ��l$ {��e��"%�F�"Gs
[��yd3�$��g;���~tG����:�\��r��m���8����{����]�Av��z65,+�i��p_z����@VV��D�٣��l �R�5��C��DcJRې��7�L]aYX�Q'��Y:��lNA霽a���
�:
˽�1��@ƚ�N�03�Bb����)K�(��R�! U#f��G�iz!�/%��+#;t&e49=����A��*�z������3��>�(�"�u�EM�f��,�K!o��l��̶<�1[�0�-k�yf=Q��dd��g��( �v)!,���B��h's�`x���E�m푑��!N�9Όl2�N5��Հ*���#����)��:c�1��\{?T����o#'4��7iի$�>���I��K���LU&�����U�D�^6Ȃ~@����~��3��%*A�G�1�0�T�;��9pn�A�(���$�a���z��?��Aa�fj����̬p��I���[ꔷ�ܕi��sf��*A��F��>���4���}O��z��"��uB�����>��̦,	�dKdY^e�8̉;@Ra�q8d^�����q��nT�2M��R;7�]�`�Ì�8GC0�e�ei;gߞ��r��Ʌ�� سЂ��3��_�ئ�fUJ
�ͪ	�_V>�� K�Vg��2�mku��?��cC�h��62���j��0�I�یeue���E7��7�<.x�{�Wn��'n���~���{�u�K��'���'[�6���p���No�k���0��S>���,�v�5ٙB�c ��\I���CL��W�_����2F9H7h=�g4 �H�0����i%��~j��$��-!{0#�&r^�L�=ѿo$ �����YV��|8��؅�4@IXl��6u�\�,f� w�YFN�r��g����.cyJ5���A�>�����,5�x݅�� [hj(�[�F�w�Պ�1KCz�5A0���]Ru�9�b��FS���~괚��Ҍ2���k��Hd7:��[�t"pz���YZ���n���E0�%�D�}˄���R�9e�9�l F�:-�Dd���ν2�g�Y�g��h�Cd�
��a���a`2�\1�� Q�>�]`�DT[<qlZ�+`��$-��X��������y�Ey�8�� ���I	`B{��܄N�[u!t٭e���9�b��� i��.�2q>X���&{ݱS���'>��N��!t��W�g��N�{՞2��S� �F�W�d��dvne9���� ��+�&o��RQ�:��y����{�Θ��V=q���ר�g�ꐵDy|iyQ���{�N9����@`B[�0�74 %���ӱ�o���r[�A�?|���x���x\��G7n�����w�q�j'�?��]hO:c`T�>U�P6��f't���ٶ���Ơ�ӌ+���<&z�F�o���z�a���C6�_�<�������s��*0���K��!9�$A��,WX�<�=�^�8�ss���9ba C��!/�ÍM\~^���M����(�|���y�HjD�z�W��`�2S����ʿzst#c��)u�)ڐ�{煍�v�dT朜����y�^�}^.��z"匦�;�&9�
�l��:;�'g2��?��Q�q�J��s�feJ���,�z.cs�!I)��j�&���pC�������5�]���y�~��3gI���e5q�E+=ۓc���P��3����&���;Ή��gY��
����wc3�K���y1��8K��8}��@`�?�|�B���1��ݞ�V({��ܳS����ܲ�k ��	�N�˃rd��Vnlwn��4�q�s��wy�Rrn?ՆLK����G@\�o�!����'ZQz^O<�V^�F���>� *����j�K���=�si�d%�1�Ϊ��x��wr���]w�=��������/yF@卭�LF�� [	|��3kqN'��(�R�5��:F_��N��1�l�Pڝ����bN35�{x�rZi�f��C��N?gY���=�rp^aF�(�}ߡ(�2{e�S��?o���(����P�$�:�u�3����7I�)�A�^� y�����(��Qڤn1�?��ê��n1e)j��B��
���UC�f����z���^�s�����ū�yY����)9�_�d}�Q�Ѽ��QXhhe�y)�*<;_�A�J�v[�3�^C�{ޔ�t���Zx��2�
�V����*�9����x֗+�}'+������=�$Q��ln�f���@r�^"��>/�W8� A�Xf[E�#�a�l|Ԣ�;p��LJ8�7�I���=K��Q>#R����gFs*����>�g8�bZЙ؞Ꮆ`	���J�Y��C"��z�\_@��	����v��=a��A�;2�Tmqk���l
؂�<�Zv;���I����֤ړ��$�8wmu��=�s擔T�Q=����c<�*�q~�Ɏb�@��b�X:��67���$��}��x�s����/ߔ���x�qճ���O~�3������.���(�%.�d))��`Z�>���3���`�0��Ӡvm����Aco���E���<
��o�Y���dş��i�(߲�³e�ˉ|����?��ܺe���g,SY6��~i�oD�ee�ҹ;�n8��y>��Ν����V��*P�q?����]6_����J��e��d���-#��.�����3=�3�r^9�H��C@y�Md��]���݊R��VH�ϱ(\Vl�O_��K=������ys������0.��<��R�#w��sg�*G��~�����W� +1�6W���lp��%��Yu�+Q�U0Ŋ�Wq!��ܛ�(���ݾ%QH��Q�rfχ������Z:�¯�"K�9����Rl���L^12O��1F1�;���6� ��' ̲r�`�r��K��������Xp4�C
�H����Oa3�l��-~�נ�3���E�@㔻�unh���ƬO\T��=e��|�l�3i5���
S�2V�R���<�"$y��]��5�aN�e�@N]u�X\����ߑ����+�>.:^w�|�M���[���νh���E���`��ȴ0���{��X�"l��j>$����Q�����0\C��	F�@�W���tse�y^�.��.�/���~m|Ґ�~QV>���b�.��B����Q���L�v�<���7��2K��eZP��{�[�Ye	�e���u3�0�R�oh�}�벉�(3z�@maL���J1F�.S�Ls�M��eaT��\��'��ݓb&)��Qq�!s{��Xf#E�S,G;P�(ת(��b���(���.3���.�������9}�9 �Ci	�C���dS���4��s��C�.�*H�$v�y��^��q���!tc�*�H� ߭'Wn�i:!P��w���*H��������:�ѡ�w{��=�BJ���2�s�%q�?W�(��
OTTȴ� ����t�V,�Ǚv�9f�����+�s}|� 9�\��v��E;��6Aͦ�Jb�(p�W�D�����@��n�(G�b�� cy��6G{�R�@/��7�T�K��d&��O�s��]����رc<'$���I�B����&7�bJ��l�����lwaU.���;�~�e������={�88�1���g��rQ��-� yGD�ɦ��~�1P�YH�zA�|��H�F����q��ƕ�/��_����AF�����G�*dΐ��Y��r�);*:)�
���
��򌡧$�%��3C��#�3��YDC�Y���Y��yU^��=M�s����Xeӣ�)����5;���ЀD��)�1�b\�E�E�Ww����ʉWT}�y'�Y�㜭�����J�e����2G4R8Jǒh�~o&���>�2����q����%�O�YVGU��� �EQ�Uy�m���z�  ��IDAT%����\v<�������\y>�k��i���TS e ��U8.����6�l��\�\�]nFRq΁-��=�UʶK����E��#$Ș���C2���5��<�����BA�V�73�q_##��I���ρ���a�M�=���t�5:*��V~ #@ܿY-Gr��D�Z�R�[d�t���`�Y"ά�Pr?��ZR�y�Z�T�5�w{�J�ϱS�5&HRR� $�K)�v:�����U����D%�tL��)�0&�טj�+pÃ�jkgO�����{A����z\s�5����?��w�}�{���JY\X���m��3U�a�9�^I�������	�OY}Uh� �Z�Fq8�<N�����ѧ���e �ӿ�5����KY�+��=���k1�S���Y�_eeR8T��g�*��F&f'k�?�H�^�&�I�h����s.���yV}��ܒh�L̝1��������~5G+�c3<\�xJ�E�׳,AE4�E�3 at��n= pE��O�,3�r�ś�x�x�b�_l�H �#˾�#+3��s��`��o���g��h�ع���fߡ�m�C� ͷ3أ� e�Ue���qw�;什�e���;�9�zB��2c�J��z�9�����$u���(p��Q-��m�����[b�m�c�5�Uov��9��Q�mk�X�,;D+�]�Z��fы��Oe�y:6�'���e�y���m:~ �9�>N��;5Ǉ��_�x��_2�#�M��3-�*~J�j�\`(MIj�sլ6����s�܀� �����ƙ���ӍX�'�� �yn f�kj� .��ݒ���XB
1��O_R�@����)��n��Wo�/��z�����;e��Y�7M�de��$��x�#՞n�вD+U�2� b��z�a=�1F��f�l�}����ʃ�8�<���rFO�tx~dD��U"'KTf��S���1��>Ӎ��?�O��!ՠ H��q�a�o��gN��W��SϽ:'�	fY��[�0��Jn♱*_���H�w.����zA1�,�#����u�HP�=A������љ��=;�zD[�	�`3�yyoq?]�3�N-צZ++#��R�l��� �}P?�fS�=���ue��xv����F`��;/�.ISp�3?���oE~E&aI��>#�}�͛�y��Nٞ���<��+,k.{Ķ7l=����2��v��Oթ%��%��m���l��}�e��w�~h�擌��/,`�dS{	���@�z�l��l~�7��GcUY���'��^����Ԁ,5j�b�&s՝��.F�Цj�=E������v�YE��$�k%n t\���:�K�;�R�����@���.�Q����9���v���)���hw A�'p�c�����48g�5xP��������PZk�;�s�����x��8r��O>���9r,�5�9����(#I���0�����F��dL��zC�T4��D:(��ΖF�]���v��PM��ey��eY����2������ɖ��Oy_�*_fU�T���|�D3�y��TiQ���>�ޔF��/�19%����5��XY��A��9?9��6>��w L�\gwfF�Y�T?/A3�
�c�֙��G�Ȋ�;/�K��Rz=M&�ˁ6���ȌƩ�D�-vF�4�p�|O�D����u+s*C����Og��� ˵�w�֋ˍ"��zѸ'�������A0�h�_U�����D�j ��9.|RTR�N����~?M�9�[�V]U��h#������AT��Dv �T�r<ʐ��zu����7�α�=̵$�0�y|�2�9�rO�X��}˺I��(2�J�M����#?��-zu�h�[�9-���M{���l��g=V�Y�۾��8��M���d�f�I�"�=$�?���}�I���$Y)
����6��k,��G��_{�1i�����yM�,H��	2T��"d�7���{�ը��P�Ig!����\�U0��b�%���,v�i���u�uO���k���� �b�
9�6b����/6��EA �\Tv���/}�K?�G��uc�nyqI�=5;}jJƎ�f�'���s`o U�	Ӣ��Y!TrB�e ��h�\�p���;+���\�+�RLf��U�Ӂ(lp�H�Y@sY��@&~�QzFLPf}Π��'Sf>�m@����9M��8˗�f��i >�3�iح�[��0���R5C�zx���߳�X6�gVR�o��kl�i�mN���h���N8:�C5b����`"��6��4��j��%|n���,����'Kښ�E��~�߁Q\�u8s(�����?��N��Yf���%&;��0�4�.�(�����
� ���:�qY�50R����a��$g`�J2Ω{��W�de�yn�<�ys�Aa#i�ʬNd<����F�'��-@� �D�X���=���!+޿7��
Ǎ�엳�Cq�_E�X?�ٳ�.�*�Q\KɤV6��V�Q#u�p�u���E�����L��ԕ�JW����������{�%�(�qǝ_�e��Y�:¬+�g���J��&P!n����'�˟)_u�5���epv�>�7�(���hA�u�����믗��KS��h�IX���]@W�6��h��]|��v g���n�v�m�,�E��Lt��ҟ�U���k
:rh��Z����;6���$Ĉ;3׎�I�~������K�����fu��3�;���ۣD`�$�"��Uɧ0BS)qą3^idz�h}L�#2�	��%뀵���L]��j�5[�g%����<�<��́��(�c��\�{����sr}.h��)�o�H�N�e�j�B�J��XMX O5��d�>.����7�Q6�,~��,�pb��D��}Ą�S��I�4��qc *�a����X���A8��9#Y����ׂB���\C���Z��J����8
Eq�	�7q�!��/��Ը��^đ�x�Q�e���|�U����|��<D���X�0����P���� �I0�0~a�8�f����MC/����'#�`�N#��N�{�U�kϜ֔`���L������`�ZCsY2���%��<�k!�������VL�Z��t�0hÚ�I��L˽V)�h��D���@/��+��k�*F�}����2:ދ��3@S(371dү���|���ܞ}ɥrdmM��|̮x��PUhՕZ�X�\�|��$nY`�#'��^���_��?q��t�Y2�i@�e����x.�����o}�-�t�O}�3�o}?�WU��Q?V3����o�?q�W�����Q��
Vؤ�֫lw �9JQ��n��L�1�0J�6|��gԣ��7%,�8
���;.:���e7<|�������o��-k�7Ј3��ş�7څ��%���D�Sd���M�G�F�Yo��f�0�3t��"�+ź�Y��A	]߈����]��b��r'C7+\#��]&N�`:W�s4�iR��ٛt�S���6'��,�s��$x�k�L�~��S�+�\S3��s�?�����ڟ������W�4f���⠡�rZf8�w�ѐc��h�E	׌l��djN17��i�-/b��	L��ۋKv���������VD-.2���1f��{\M��J�Q��j:���I����!e�9�Ǉ�+l�Ӿg���k���s�����y�Ĉ �tZ����qISz}�-��D&�\F7�?���Y����뵦�D`�2?@a@
�eT�\��}��m�t��!�-xE�����3'������No�LP�l�=� D2��J���p2��Kb ˋr�+n��z�|�����l:8+0�P��Ŝ$���>S��f�Ìt��nG�֗�[n��=,���㲲�h��}�@��V�%q�e�&]�o��o�3g��m�ݦ���[[�c#j���ԗ��6֨��[닗N��2Ynԝ0Dx&S�}��g���N��rTYqܦ�f���=p���!�b�mҢ���v��{�x�㦯�����G>��e	nұl<rZ����R���N�K���|�9���ʔ`tB����d����.�̍��D*&i� r���������F��U���ƾ?3J�r�@����?ʦf�WI[XT��FȬ�����,��`�0�"�]��)�Y��
O3�q�8���5�I��X8�3��~��*2��T����Q���(��|vß�}�B�l��2��i�:���WQ�(_Gɻ܂��Dc`� t����`
&\Ʃ��${��R�83�&���g������r�����ʵ��j>%aU��;�(�"L�}�u&Ƥ��J����,j��sF�@�K܊%�8�V&'U�ó�
�05�eՇ�`��_D�f�ӌ�qj��q�b�`��"�G���	�9c��G��:��| :[�2�3���vK$�=U��J	
��$�L_(���D�o�n#��w�e�~�����𫮗�֞��ϾC�zu}@gӁ�)�Ñ, h+��5!p*�p{�+K˫�7�I>����f͇� LQ�:m�9SVg�$֠ϋk�}�<�Ѓ��������ԣ��2/��k��Y1r�.�UMP��KPu���)�x��ލ�;��Yn-ҮS|f���h�:5�S��(�t��<��}:3�{��l���r��?sؿ�����3{;r��?'�ӏ� (2�\+�3w=O�=�W!�����@֕�� ��Q���#� �6Kg��9��qE�+��.�����2Zz>��(OsN �|)��~!y�r1(}GFB/�\�L�	8JPS�L4-4#�v�._�u���W<[R����L6q_V���s����ߗ?�5�\Q�v���!W9&�������rҲ��8:Ð9C@ c��'I�����E�ǼF�$�nеN��i��(��vu��8�CZ���ey#���&FD�bO��$���C��.��1��*�	N`u���sߣ�4* �~��Y���E��ɕ��.Q\�4@�z�R�)K�X���O�8��!�g��ʚL�u� �y���Q�� .dP�$n�equU.������s�ao����?����3�`��c��c�h�^0�C��].t��
��K��Zߜ2z��`$���ߔ�C? �^�L"�����mrX�)Fbp�z;�u8�t�����\e	a *I��7��o�G}D~�w~��=�Tת�9��B9|�t5����w|������|�C��* н���R � �(�`M2��31cK�#�`P�-f���g��D �L�a`����1�1c���> /��\^�>1ޏ� ���lEP�j�E0O�QJB�u�]t���н��5��]�%�j�4���  F��n|�d��{eI�"�jF��J��u'��"�(�g��p<�d��Y� ��'f��4��]Ȥl�ȑ!�#
ۗ��%.+��^B����0 P�m%X}Ȣ�e\��Y�m�Y�Q��S���a��ѱ���6K�r��)� 
�VgFS4��F=�8������fX]��w�iitg������Z5:¿	�,��T�"W2ͨ�k�624uq�NMG5�����@���Z�E�i-,:zg�,p�@m�a/��B	�"���"���"��l�ê��B�Yϭtᬊ1�1e��U�#�Hu�X�M�zΏ~5��ң� T3˙�+��O�����=zT�5[?�G�����(�U�+˴e��u:�8�?�}j:��k����j�޿O��_�{�Ov�{���&����5�Y�y�&�h�?��X)ޞ)�w�6W��#�\��VE����= tA` #(XV`�d�B�7%PG�����>�`O�����)v��Z�a���IR����s4�C\���,��ɫ����Ï�o��~����4�h�9e�=�j�����th�;{��W�d������Wj���aGV�]I�c{P<�4���[��?#�����ˍ�*QJ� �F��%f!'ZzW�b<|<!e%�.���"uyZ�=;ɓ���9I}�M��Aҋ=ދ�?}���'���@ �հ��83A�L���H0L�=g摖y�d�.*� W``�~�A�#���E�#&F�F�7�yD�p�a9�.�4}iv:�lkydeLW.�빡t��5���ˠ�ӇS,��K��d~6!��K�,R��eޕ�M���X�EC�iZ�,U!���:�z}E3�-'}]��$aNc��5i6jd�����O��S� �F��Q�J�Š~��׎kB�%n8O����8`��@_��\��w�#�}�9vTt���+&��4���us�(�����}L�{�f;���x�h6Җ���o�����b,=��� ��mUʇ?!"y*O�~L��	-�QE�u��2���F0�k����3���P+�'�����HӠ��!d�G]p�T+�N�)KKVR���c�BI6��H�&q���Z�4��2p��'Ƙ�vR���������}���|��F��4������|�O>*�z���,�o������Iu��Rf\�Orc~�#_c?���*c�8��!S�L� =�D�A�/��s�j�]����2V���|qiɀg���XY����ż�Q�nBɚ��bs�2�(��ri�by��ߨ��P~�n� G��BC��P�)�#]������x��tu�W��."��x��#�@� �cyy��O+�[�pd-�M��lt��mf;$EiJ�k<Ϭ<y6�nHp�=x8c8f�H|�I�4>g�^l�GA%II8��;���f�U����z�n�-�n�iNO��9.:�� ^I-p�~�ץ1ܕ��Ӏ�&�L��F	ܫ�˽�	Q!z��5���=�`K7��+�9J�0�qy���h	"f,4k��z�k���LL���޶���1(�\d�俒��� ���Z|Yҿ����it�踣Y6���P'j���u#d
�t��^� �F�[jH�Db�n�p���/IT�Js�&C}��\�b�)�ͳ�?�S9��f<���F�7������_����A6�N���k��_|ܘ�|s̸&d����Dn|�Ke��1:�t��n�59�F�_����+�:y _������ч4Siʁد��3���~ӷ|�<������R���k��n1#�
�J�������H�Nl;fQp�<���u5�q���}��S#�{�];n����#XM�d�g���_�My�O�� ;��r��F_#Hu:τ�u�����	�?��+Ca3M�k�3�h���~?4f1�	�ܣT���m�.-�4��������ў�k�0�>����z/"�Ud�8,p�\z���Ⱦ���/
��6�C��u�'��a͎��%��9u���L��k`�'��uQS��[���mr�]� ׿�i��Q�D�>r�Ü[mu����a9u�eƲ��i8�P{,w~���?��cuuf/x����� �#kz)cY��Ӻ�V5���?�C��:��m?&�nK���r���t�\���?�����Ç�4�y�=���Q1@{����G��^H��z�5�w1��.����f��ّ�x��j�Aq��pK�Y�6G|Vڍ�����@�U��M����]��ృ$��2��9`|�]�W�ʡ�"u4�4��9�S��o��A�kd�"�q�s+���24�7 b�jK�x��ZV� �fa�_�{���� �L��	p@O��ɢ-+��k�gj&7wwj@9�'�q���3G�G�͈j榡$�3u�z����9��IF������Q�	�ptS6bA��� ���=u  u`�Qr�<����WĆo������F<8o�r���^Ї���
�z��k�nU8i�����Tg���.�nW��9��IZ��_�J�R��J�f�� %*d�����:�z�ô/�!BK߿�q�@?�5�Y�4c<yN~�?��V�W~���Y^`������������W}��8x�k���:g���~H�V��p8��3���m���w���o�Q�k	g{Q�\�5$j��<�/�G�����W�o_�F����f�[��_���K�$ߕ}��@?�I�l��l�:#��^�>u.�|�7������^�^`*3��t�����-��	25��	ztM�RǶ��jY�&� eY��P����M��OlL��U����iֽ�f��}Dvu/TG�J�f��@��W���L{F����$���s�=u�<t�]XĲ��q�G��Y����?��e��K�����ˡK�Q���������9�]!?��w����'k���|�����"�V��,�>��
�{rngC��-˫t�k.�D�d�Ց,���ǎ��C��8Gr龓�J��o�_��S�Nɮf�>��<�W˿����{z]������w�������d��4t�~���ʒ
_u�_�ߌ䁿�C���_�gŗ�~���ҡ���mK_��_��wɛ��Mr����ht$��ߑ_z�<v�I9���}n��I�'�;ĵ�	���l������x=��z�k�ޣ�k��k;�2ل���xW�^����_�������W��:A8t"t�b��>))]�\��Y�x���`����p��x���x�f�QI�������A��dQ�0hʌy�Ҕ�G�%����y��娒~�JԒ�s{j�����|�t��'X������tG�~�o[Xd���<�)�P���>����+�Ob'����{d����R�1�A���{R��L��c5
`�aI2�����c��t<d_��Qu��-(3�C��X	J�j�0�[#��v�X�#�������ͶZ��x�["萔e�T/mO3�Y�zW��C^���1�D�z(+����;r���_�u��YWț5h�-���i�{��׷J>�����~��/7.g]���<�YWj�5�I�ٸ����s���>��w�S��3r˷�K}Jƃ� lj"��O��_�
��[^�k=�v7IҀ2�+_w�f�S��?�Ky�Kn�����ވ@���mK��6=��%M5�}?��SZ�;M%N9S�@�&����-���;��^��TS������Iٿ��k���OJ�=��ş�79�q�\y�$e2R���[W6�<C	Jd�yݷ���d�Ҷ6�۷ʿ���h�p߃ȓg�������7�A=B*�о�?���/.�ZwE677�/�ǟț�����3�K]��ÿ��r��/�g��B�z������}���%7�(W]u��s���_~��F����5����ş�y�s�+_�ʯ���wR����|�O���Pg|�yW���R�Z�h=�
��|�_��:�%�� �2@�u��W���z!���9����Ӻ~�-?*ϻ��A��{�w���������7�NoS>�G�/?���<�yϓ��M3�uz��?�g��:i,td�N��D��O��\v�Y}"��ٟ��5{ٍ/a�7�F���y���O�]���?�V�>�-u�#�c}DJs�,�Ƣ��zͦu�.��~�+���;��OJW�0�&��Pj��w�N1��$Ҡ���My��{y���C2RG�m]��)Q�2�m��E�
5\��BD�u!�$D9��*��8}͒f�p�,W��X{	�B�(h�����g>k��C��pL��<d��z�^β5�8;TI
�v#qP�=vo��#�@�����9�k(١�J"�xHͻ2����ӂ=%8I(ǀd��kB���-}�:����T�2Їfk2�^��X��)��جk>���D��7�y�2!{8��f5�-AÇ(wm�+#������o��D5�%�s�,��n�æ�m+��f�}ϑ~������X�V��4g=�1 fj�Qbm���K0S�g4`sf{���o>�I���������H��,,�7���r�=��C��G�])Ya_`����^�H���}�<�9W���-]���������L`����P���2��s�3�h�׵�����(?�o~@�����k_�"����qj!�É��.�I����2!*��#YY^��S3BdzK�T���+�ӏ����M|��>y���}P���?!�r��q9�����?_N��zIj��6v�����o�w?�u��m�w�؏�[~��r���5��������s�o�.u���}��?�S����M�ɟ~��ܽ�G~Xn��������o�d�|@��K�\����WM��$����$o~��军_�s~ε�� �2��=�k��\�M"Xc� ���7��+�` zr}]Nk���D~���d�Xz��}`?v":�{�G�j����Z��>�z�I'rN�Ƿ��;��ӧee���y�	y�{�+߫�~͋n���])t���8)����?�?*/��zYV��η��@�QoOF�;�>NV�K/����Dǡ�,��������뽹�� ?�#oU�'��X�@��k0�{q�חH�ݚ�ö:V����8�:���4P��5�LpCFXKu2_�қdU�O��t6�@�+���g�< � �4vk{C����d��qy����ۇ���T� �[�ƥJ�[P3�)�*����'��ي��C���}VA���{�' n贝� h�����Tl2�; 9Z9ϱ݅�L�cC�l�+G� �@��H�%jwX9���d�4����x��#�R_7���)��
 M�n���U��M_��h#�*R���/ 
�{YB��@.A֧�2U�� ��*����f��{�ᡲ���f���uBat����YQ�����~(�0���Ɛ���Ld�a����.-v%�M���9}`������}.�F��`�態�G����c�=�$;�k�}ﭜC�0=9�(��"
H�@$���d���y`xaLp �1IH	�B9����=3���rݺu��ϭ��ߓ߿����>��t��u��>�9{��ͤ_���R�pc�}x�>\�⋑�M�F`�2��GR���%(�}�_�ʥ""1P�,z�3ڷ��e�UZ�B5����vaA/}�ˑ��r] W&�D&�lt~��pe��F�QJ��{�VVg�	�|Q���V,Á�q�%iz�
궊�0�*�#Z��o7~����jQ�[_ s���k���a��tݛ���9睋��ڊw
HZ1r�N;��B�m:��z0���?�1.8k�}��5� �x�+_���)l���x�i'�b0ۋW\q%N�	{"7�x<�K^�Re�͚�IKF��_ߏm�6�_�ip����oVn`�Y�Z����(y�yϯ�p�E�aکX�|6�x�J=[�����zO�?i=��^�ö�N�E�m Y� �U�u�������w4S载Y���t\�W�����2����}{���V�#"�?3�#�1Y���'����Oـ�o�C�,�ͣ0�?~��8thq�N�PL�qx��sr�1 � l�0?]Bvx@��:�׿�J^�Ρh\�-C��"�\��a�1���P�m�vn�y M Rф�hK�i�lW��U��eD��in�zI�\nq�g�B_��2^�Wc`�|��C��)y}M/(�O���[��<Tcm	ԌY:��V>_�#-�홏,�:��2�gq[G#�*`A�C��{@�+E͸�Y��`�%��v��:�6����{�i�]�\� P���gճ�cD�I]�S�{^��q�J�헽�-�q��.��0lS�[M�^�=�T�T#����$;���F{LK�0�ik&���VBAn��dF��|F$��0�� u�QC�Q�Dߎ��Pp�[W5�Y����L/��b�l�V���=�\;�Ip�'�a����Ƣz,LC����s��`er[�8�cA�C}���^�S�F�]�k�`��w��|�a4]}m+����+�ۣ�x��)A�c�d�r|�w= l�tN���6\{���t�U�f���~70J�ÿ}Hӛ/��2e�f�7����h�vXXTO�ퟷ�^�M@���j
�>�%�X�j�:���LO	b�W,�*nϐO���(��)�HT΁�옪B�RZoH�۟�����|߼�+8�ҋ�I�-�
 �X�n���҂w��$�!��{��	`М�T����0�d�L�9��Yi�D���C����q/�a�/���^��~p+�����(pL@k��U��W <ԣ�U{>ի����;�rW'�~J'�Uଠ�T�ZD�֠f[K:aR�l"�X2�K/\��7jZ�U����/tl�R�V���Ԋ~yMv�[�l�?~�s���7`J��P۸,��cmhA���jr߳r]"[|��Go�ox��]�����������k���gl��s�<2�+�9���L��� v�م�[6c�V����)H �����]��G��zE���c�-ޓ1۫��N!>���EV���F��,.��
��af�EI����Vj��S��@ �4E3$pbA&(Z��&U�a;�i�Ҝ��0X|�����ܪ0�Vӫ�g���1�Dh��Ǧ�3֛���L�Q�/h�������9��C̟=;F�%��7=̖Z#��S�����my[�	1�������S8�������wv�É:���ñ�m؇W2O�I�e��I�w�=��.�zR�
:x"	\���[4�v��
��I�,�2N�G�Fk�{�l->��/Ӫ*�Ϣ���=�������u��#�u��Ý�GJ�̀�/�5���Q�ʷdⰽV2vyO�\Ԣ��LR���s�^q�����������>���}:0Hu�Y��B�I� �j�H(����_��	�e��	 �Z<���?�)�n
;�	k�����l�!�1u-��󲫮��SN���ʄZ��5m�X��`�%F��r)��2��Ja'a���)�  �g�֬;I&�(������,r�19΢\��/��Y��0���\X�ip�u-��kN:E��4<|��8����Z�Ut�B9�@T>�S�å�h �,�jW�r��5�_�ª/�r���q���{>�?������O']��O�H�oto{�;���Ž���͏��}���>��ϫ�o"����������RP�8� �gK�H�.�!7��ɵ�j֐�Ia.����n�����^�K�'�%���\sC��/,����y�h�ZQ*���}��G��G��O`��5���˳�W{���#j.B������{����L_z���j�X&�\� �s%|r�#����S�3��[-c�)��$���0�r�6��cLw���K\���:.���.�k��E�Y.��"�ȹ;��i����+R��IPdԩ.�;H��`{KH�L뷜�(����.#����sڙ�BIS��)�q��a �Xq,�[�Br^��������ͨ>�uܙ�].a��v
��Ь�f6���L�s�rlzE���v�|�U��O�Jvz�ev`�J���:�#!�z�d���2��۸�=�����o~
'������͎URR�}F����U{6`F��ӳ�z�����Lo��`ݖ<0��Y�e{Fi�ܤqNVH�����$�50��CզD�m�PS�)��k�k���sK{4s� ���a��%���Т"M3�@GP�K�o̎��lC&΅�%��ͣ��-���U����yp�@���i�Pc�u[���;L�OONa���([Nd�d����d2�!��̶'�Ľ�I b���ڕ+�f�j���ߏ�L�u�LȤ�vPeц	S�3�>	2"
b���"p6��	�����Nbh�_3`5 �4��<���x�$�d�:��;�M�JT�D峪r�(��I�Nv�3o��9Yc��{v���{w! ���?�[֯�,��z��t&�k�a)�0��/y�8���.�z�����<�	��"S����/�R"��P�����*(:4. 0�����/�b�m>��)�����my,���[p��oS��@ ��#a�N3rE��j{���J55�pU�!- qdf
��������M���= ����j����N&8_������/���sT�%�w�+��m�ܪ}�gl:]���CGp�=��uo�F���E"��ܣ���lظ^��;�|
_��?��5w�7(W���M�=�l�Fg��Uo|#��կ��'��5�}�
�}��0#�b= �"%���^o>A�~�=�������E�c�� >��1,C����T0ӊa��%�hV�h�j,ڴ_���bY�5�&L��;ecr�zĚf�4�az�\ˮjM�fG�@�y���޼�6���^�J0�gJ�ٖeq'�b�f��/�<iZ��A�Q�;*Ik�m�kO�R��܎[[�!P���ذ�r�^�g�ٔ{���P��낫^����oq"�.������`f�VhQK�JF��ou=��c$�['9Vw��ǫ�˦'�h	�Ζ
Z4��E����Y���~���i��Y���	���Ɨt��y���T���G5m�@�X%#�|o&��+u���D�x*ג��@�g=�̈����R��(-(,������L����,�h�Q�ϗ�4)��5E&�/~����I#�J̏�L$NޠVfq�9afM�I�Ӑϝ��1&Alh�Fe���4|>]�Ղ��O�UZ��Īk[	Ơ�EV��r׽w�
�\c2�%�&{T%),��w�LN�ɧn@-��9�����P˔��E:,2���t��W�N�����~WC�>I�\/�_�.|��x�K^�?����;?����W�&ݭ4K�{�A�3���݊իW��F0�BQ�����fq�{ޥ׍�r�J	k �V5z�2s!�(��m��=��
����
ZP1�T^֜@�?KX`��'eQ>�od�\�b|�_P=�E�������.����/Ӣ#��w*�D܋3���H��0X� "�M��tN�"	-	�jXu�r����O�����e˖iF ��-�~;B}��8��i�7��M��߾�k�%	j�ڲ]�2��&�-���x������'���}�߄_���Y��%	"N=�,5U��^ϭ#�K�w�?��V|�G?�@(��]�:�⚫5�P�fq�.�!�}�$@���ˀ����Y�^��a|�cF��"�"{W�R�i��ӵ"6^p6��ی�|��K�1 �HB��KC*2��L	h�Z�h;��+�9i��QeL�y&��v�7�*cf"���V)�DgF��_[�ѿ�K�,�Q�4�k�650L�ҙ��r�H��F�!��~p�iz����V��m��I� ���ܳ����W\�g6�|t���e���2�V[���MmYUv�B�s����&p�j�Ƕ���!��	���ziM��|�[�a�M��B�<��rE��znA{m����`�y��-7��ʕ���C�M��=rYa�	38>~Pې\�!�����L��[�db@&.aT��+�ˇ�)3
�T�e�t��f�g���8�71ӥ*k�3����_�/}�3X�d%.�+�p�w�BS��J����İP�[HS�U����1;7�83�P��m��j%����*Œ6��	���Q��߉���_Ogp�L�K�1;3#�_�-[�o݊7^̘�E�*� ��l_�}����Vd����3X-�P�i`�PV����n��.`�I�Q��f�0�H<����JL���w���ߢ�(�8}�22������P��_�~���aÆ�V�u띘/�q���b�ikP���t:&Q�@������?܃�_s�~�x������0%����ַ�t��X�2�%�l��4����k��W��U�N� �L��z9ξ�<�\F�{+��b���t��*f"�Z�q#�^����&gU�KV�@�)0����/EDb��tY�zzq��g�gd������˯x9.��b-�bk���5�Qd���ĕr�?��c���J���u�����fA�M��׽�-�؄����Q��R��3��+_�j�YP�5����qI�"��cHP�s�I��3��$�����;nA�<'9���4����,���3���λ�r����;�x���G�Y�I�J��Ug�b<ͶRYӓ��`���2��������]k�{�溮7��%�o��
g�q�qT��3ڪ�
�P��
KͶq����т�E��^�뚰+�%����c���lŹ��DU�������V�[Ϲ�h�魭�!q�p�c�f[W�l�����<��nS�'C��4J6� ,�i�c ӣ)[2l�YZ���s���#S֪�d��#MWSǮs��n�:�!S��[짫a^�4�r)�td�B�O��Hm����esߩ]E���>�LS�'ʵ�`L�[\�	��7����	}�̰L�[& 4ZO�m�66m�m�6�m�f��vO���l[�}���|a��g����ZN巹�i�;����{'���z�үĩ#|WSr�|�I(���/�_�MD�Òr�9�Q�<y��l!N��������P04��?��-'}0�%�B%�q�vr�����[F_���3�^�>��M*D{d'��ײ8��ja�ԉK�4_�a�X~������V�,ܫ|e\�Qh�r^������V�m�w�SA�Op}���c�f_��Z�Kl�3��=�\����}"�0���վ@�^+}��oA	36�vxYчr��DMT��3]�(�$"۽ќސ������y��y�oY�w��X��[v���<�l���>C�*�G��È���S��I-�%G�5�;����5�09#��ͶE�e�!`0%�Z�T�+Yч��N��DyGx���p�ِ?��]��JmR��OC� ��r:ʄ;��$0�������5��e����*O�����k���&�, 1��!MF*7)���	�p��	�������$�����iT����U-b2Bף����(V]*��2��[R�־�SFC�~$%!��頳�|!�3�O#��p2 �j�ѭ�\N�� �`ݭ��K�x���������A�>FT獍g��4h�)�ߜ1�Ֆ֑=��g}�1�yw�k/�}"G�%-d��T�B0�j���
a���3��s��Z!8.؁�z�_<4�/��ȧ9?9�l�?�;e���*֖�����\B'��{�վjVa�$����L�To�oJM��@.�D�u�k�s������J|�@����KI��*ވS6ט�N�
o(U��VؠT7>.�BF}��'\��[J�<3�,�
�MO�i�f#~���M<���E�ǤeL���;T�Z"��&�hx.�t���eN�@���������#˜�j��Ϛ�.G������YQ@�cv
��!���t�B�97�	׊&�i��aՋ�oTXD�y%xi:؁�����8���}W����P�גF}p�HL��QRp�l=ϊ*ܺ~F���x��?��x��?jB�P���ٓf��!���8��WT�Z����bP6�=�1 +��<�u;R!gV=�>!�����*3��ztp��鵽[��\uJ�Q�r)��TE�Xa�F�0��%B��t>H^�,�m#�S��	2,k8���( �O�~x_r��8�/H������O��/X�>���>�0j�(`�I����p������,0��ˢz�5u�h���j���<`�TG�8�/�^5�^���h����y�UCl������u���5��O]N;�6�}�fҌٵSv�a�K�ĚY�ȶ�����#��O��8E�޷�ws���֓w��Lҋ���jBg�̽�<"N=:�]�гb�M�2��R���Os��yzCz�	����-�k�C�=�
J?tk�O ��xZѻw���3բؿ��u�i'ru�L8�M���A]z����n4Xu]�Ӟ�P4!�H5u͗	������)������\#a}�܇='�� �ߒ��{1o�vq�+Q�{#\�>Y�~���:��7l�:]$��!�}��� ж�)�R>.�a����g�s4O�q�����Vpc?��X����=Ro���(q�rH$�gi�xxl[$�"�&	z��ilJ�K̹����ǟ{�;�X�vڲ��`M�V�K�0L{~_�J��Mui47��*�o�ݳ6�* ����?<[{i�-K���3����l���B��g;2��A!d���I�w+�"n���V��܊S�H^��F.�\K8��6��
�܈u�h�[kUHYB�sS�����N�Gj<�z���'^��"�K!FM61��楅(6m�$U?Ʃ�'xbt�ʿ�ɵhN$>�?)l��U�Ԫ g.��9	 ip�^�hK��`c��M�L-�
�� �Iѐk*8W���,�S}9]}��,n��m`�O��dÁ��k�[�>���\��+�(�$Y�����v6�ȵz4:k*j��m���JmA�E���-a�u�o�Ai���P{��\��z��l�{��q��j���b�'vӑ O嬼g�4D�:|�ٟ�ū���]�\���h�^=/��6=>\�_���_�6���Pz��"���JJ�IO]�2�M1���}0��g���<K�	Ψ*A�{k�K>+�E5�w�O�
5���,qt��3aψ��u�=���͙b�H����,C�i�c��s�S���\�z�юe�=G���X�ΐ|)Fg���,J���F K G�ќ
���S�Ycd{C�	7>���ْ��/A����&N�9��ˎ*�f�����x���m=����Qui��.�����e�%�����̉�"��H�~~�0��?v>]-�̀���7��y ֓�5�CY��n�f��$��#0ƃ��N�y$_���V��L�O��_�96<`;ÎT[vR���c ���N�3�P��H@��[�&�{u=2.J�Nƶ�9��[	:��7�,�~�׋�l�2\�����,,���e�e��x����� � ��?��X�h��V��H���N��"�Ƿ\�<���3Y3���k�f���Џ}��[�e�M!"I�mt���^�4.d$��l��q�L��.��GGl���d�A欑=���%޿��U�W^>�v�=jD�y��lx�g��l&w<��0R�xrY�~6P�&݈�  �ö�rAR?q����槣�]��߃�PZ��������e)����"t�7�P��s�c����z�feo0�y��L����,�^'\�?F ��)uf���	����{�Pe�z{��ws�K�PL1��gY�cb%��\��>��	T�w%�7��Mqf���'��&t���x�/����O8���H����D�(렼@M�z�(�>�4��#�Э8��1��b���ܹM�B�����v�S�%F!Ȗ�H ����S��3�����5��tK~1~p�����1�qwf!Q�j����ong�6��}`���[����Q���쇠\���.�us�uD�g���q����#�@ȁ�FJ�8�͡�#+��d���B�|���`%����tkO�(c�	X9�+���ZJt�?����(��!�����y���\��`��b��}�î�'����+R 6�U1�PR�ZJ�Ů��r�aW�n(1���;�
W�����=[쉰�W�F�WL�����L�,����~"�:Y�H9�.܇i��c��N�O���.�m��&b��W80`�jR��
A L
1�
K&e�����N�>�1�`���~KM>G{����[�1��/C/.�^	LÂ�hM]�u-�����ґ%H�{ڲ��I���d�	�Ʈ�C�[5��(53V����x�KW0OmeyxY�M�"2y�Wo�yW����_$C�r����>�K��02q;�8�ZDf�Al����4P���D�V������b�4�e��pW��� �����_t��.ƱnJ�R _��ί��(�aBtEV�}���Y����~��D&V�<QS��|��>���g�.�&TS�a�\�����6��A��S2�ש�4^�8w��;r
D�I�[�n��%����l�F�C!��g�,��8�#&	U�>l�q�A8�vUu����֧q:깔�����m�7	1�nb]�TL�OR%�lؗo��<��i�
�[���"��(m�q8v�e������Z�ݒ�4y�x�SׇW�0��U���/�9�O��P
�aC�F��|@?�j���:KR�}�Lf���H�W���"�MP���n�������Kͫ�M�iY0�O�?/��n�rJ���,asbћ�8L����\2d��q��y��,�l<����(����g)p�v�$e�'亳�!I���z,�!��Kj/�,�A�0w�����A4�l��;0m����+�Q���~S\�Vg�-�O-E��ؖ�"V/?��a�fӣI�d!u\��(Fm�O���^�E����p%d9[n�O��B����T�ү���c'��L<�/o��~k�Q�����D�L�x�Ĵȱ��Y�H�	K+��џˋZ�SA�4_��\��*D�,BL���fV��Bc'�1�GD/|?-֬����6��M�ι��J�k�n^�&c�3gF(���1�#D�:�R��˪T����/_"�~6"�}"����MC�_%��FiN���%�J�o�]�>L<�0�Z4��:7�rĵ�O	�峈�H �9{���l�E�}ʕ�;8��c�&)����0%MVR0"�X���n�r;�&<OW1�g�&(Y9�ʍ�Ξ	��#��6�]�������<�k��r�l����nBs�u2������ؾԚ
�WY���7
F8�Z� �'�?�8mQ�o�L�����}M�k��+:B �ޟMd�ۍ�X���Jq;f�X�cm����g�K�i�Y��J����	����c$��b��k�x5.� I!�p����z�G���Yc��6?Mʓ�webdDm��s|��)���U����|���b�v>� �U��dƼ�"�E�~�RX!����WK�lDAx rk���.k5)���@h�<��c�;�m�o�
�1���\��ں�/{�]@�D���u�Ϗ鹁�6�v��jx�po�.���za?ے���֓?�1�� ;G,�by��eNB�Ӹ��0����d�v�s+A�fa��ã]8�C�)	�T��!m��pUwv�,�k.n�~�#
�N��c	?��?5�s׻�K�f��/C@ٰ�t�Lϖ��$���j��b����I+,f��y���3S����r������,���Q-����'�qѺ��A�w�C����;�v�m!,l�d���E=�x�3�&v��x�����S^�pݙׄ��x�["�ݍ�f͜��ƈre���Lr���@H�Ba�c Î2}ϭ�n�Y.�J�����[���	Q�\&_�r������ai���i�o��N��B��b^g�d�a��b)���D�fp����%��u zk4$�rY��z�j���/!ZfX��YAnڋ��|���w;(F�FV�B�j֒���Fp%��L���=u�=M�������7{C�Q8&�]ڛ;,5k���G�;�	��:���\Q�s�ocR�xٖÕj�=�N�2PBt�_Ĕ��^OkV*SǍ���|a������7���z��ak����s`�LF!��!���|��<%D���yJ��Hp�ȧ��� �tp�����⍿��<+e���E��V�R,�ɞf��X5*'{�8�����z��^�,����%����B�˪�G�c��׍v�|"�\*�,�,��(ϕ�]�^���v-����E~I���*�?΅�%��e�8Ń'˟�`��k;�+'%���lfz���y0��t�?���?/�i-
>��~���}��_Xb���u�*ܺZ@�=�T�X��Ȏ.�a�7�O#R��(F�{�GHʸ�od̯i�Ӎ����t���5���K�c��`���,�K(���x5yj�6������K���3�
�*�I瞜M��gG] �R��=��./`��B׶/D���9����x�Z�T�a'��X�&<����6Z���_���ZQ$�L��򗮮-:=����g1��1�#I���U{LL���_�hH͑h����ءJ;1|^�������dߠ�0{�^V�(�(V�V�������#�c�G��RG����CK7M�OyJHXJ����AN6�ZAv�CـJ�	|(^I��~0d��ð=T0�iL^�䭖���o��K1|c�XHaw9!o��I��9����?M��
�㏙"��h��
v���?�=���	��uV����le&d�Bt)Z&���񈧳L��4�?�ؙ����kk��,A�3�p���oP~x�S33��AMǇ����K�%�&C*�J��B�꠪�0h	Ї	5���l}|g��֗�&K��Qe�%��!
^N�`�����-j����k�Fl���s�>��#��L[~�x2W��8���a� F!�@�y��$�62Fc-�l�En�M}���T�,�a�xSL�s�	5�Pe���Q��1��w�r�ی�������$8��RC. ��"A���}��i�i��!�MN=��������9���6�4�w�~Y�F�L���=�jT��QU�w��Һ�,�8Z4���#�˘S%���T�f�}���;>��q'��/;�k~���8k���'�w������8�,%Y��UJ�9U�a0ud5����p�UvA��l=�0��>�UקW�p�f���*NpD��k�ᨚ� �������!$�Z!�ɗ$)��������~(oC�yUھO����;m|���o
��M�~'������S���`�)T[Ⱥ]�f��P�S
h(13>����Y��2�&�&s���.�ה�S0=����K�g���ઍ�G�|�I��^��x�,���I�6Ԡ��*3��9�����5�	Ϛƀ�$��Q뉺'���Z�
�(��EA��Xs����( �T(A�r�K�:����tpҢ�o�9Hh���g��n�G�&��n
�)-i
�T������ik��*(r��h��7ں�I���|��ן�R˱�����E<�}��)��<� "�Z.8vs�=�%���Km��	A�}�Vf,���5�`��6�,2��EѤ����?���9�����C��
7����3�
>�V��E["��T4�����x�N~�֗���`FQL�2#��وB�{�9����Y&@Q�7`miSڈ��f�^��As��71DDӵ�T���^g�V����5]�IƐ">8R�-�qU�[�c��l��U7��J"%\���䗋ּh�ģ,��K��7�����}ԙP`'��} >j|�il���|o��k/}��P��Z��g�����wBl�����/r�i֟7f]C}m��"�q��.@�[�|��b�
P X֛���<{����
�d���Ҭ�E��s?\���8wtc�����G�b�2��Wl���S�`=nz}L���-��Ǖ�4K��[�V�,�i�nz޸��-h���^d����nXV��i�֕[ST,����ߣg=⎛5���?�c���=l�A���z͖5P��P,gT�����E����Z���䤺�PM��_��&�ڵ���9ȑ!����K�YKp�\ޫn��M~CU���E�F0�ӽ{�f���Y\5kT��~[�N?�%(�{�a)�y�&Qc��Mʨ��IA��ϚDt(�T~V�Υ�?�E��7%�T�1x9�֕�d�(d��󮱨�����|�PS�~V�7�W
��.����$�s�aP��5#��������֨����7u���m�Ȉ��t�hݟ�?��ICEh�V�-�?�k�&+ wu&�8������r�����Ѽ�#�P]�D�y�-�&�Iƍ/�n^�>yB��B�#����W��8n4�~�{Ț⿦�9�_m2�_~nw��m}��|�
߆�b� 
�#fٝ���k�m?۽P���=Ȧ���^Gߵ���х\��d�w��g7�{�L��|��S��_$缲|=�v���wj���1������v{�w�#�	\WD=��'��S�
�a�娲)J^I��I����c�CZ��� ��H�.�$��Ӡ�hf�����n�V�B8���v�.�9Ƥ�Zvt��]k�÷o�s���&��&��[�e�lh�TC]aW k� K�8��zdz�O���@6V���?���jyq��������Pҕ�B���)��{T	��Ea��?��M��AAa��8��h�vXYA�M�&D�eBh�� �z,"p%����mTE2��_���k�Ӻ|_��Y�33����qT��[zw�ɤ���@r��X[�����)�B+O�����7^4��)X�\�Sى)�Քt:azm�������+�Y'�s����?{�
;�]
��,��-V(�z�v�
��U���\1��lԩ�n$��+��o�8f��n��)�b^sGk�����z����m�2�o��%�:-/�K��A8��;aY�ڌ$�C�U�ȼU�Ӹ��y��^?�`P֥�sF���6:K�)S�%��>�7&c��Z���)Ǖ��0������f�2��WQ
��`?�c&��TH��5)�݈�� ����Z	�̐���W����,.jE|B�[6�E"e�{��첰	]�:v^q6��5qI^pB�f�Z���a�Rr�v�0�țK/e���ћ��u�UAL�u,Xَr�=�
��
�i�^�,ǟ/������XF1~��Z�r�y��p��~{H<�΄�"�*�~��;�����F���I�XI�5��)�����Z��#�Hs���SN0-���r!_u��ɸ�8-�[ڇ�U-��Vzxv��1��oo>ƚ����s�a`��gK�V���s�xx�	+x�#�/aM����w���l�t��0�5�Y�v+���f̻�MLu���mme��+��6|F�QZu-+'R)���c֦[N����#-�=ӽ���9�4*��[N�O��ݬ�l$&~�.���n�^k�u%�Y,��+����'�-j�]6+��������L�K`��o.5MH��A�cڒ7DT0n���/��Ti'��$~��=����Y�����/����u6a�� ���@��%���cp�>�yvjiJ9��<��^��Jv\��k���~I��O�3t脮0�g�T��Z�r���{^��
<r�@}��r�۬����x_͐�}'an���y�Z�Gw����g����s����w�VP��~�2:o�|D��~f�|::�Q=�'9�Wa=N�.&�)�X�<��9��3�N,fR�3�*��B���(vv��ߩ4Ɉ(G."�x$[�?!����[&��zW $�C�t�E�3����}2�Hh��Rf؅X��A�Z�{+M���HI?$����t��Xܙ�k�N#\N��J�I���P��|�M���c��!!�9�Y�����j��ޫ{�je�ǻ��1=��X�<���7���,�ةШ~�b�Xk�LE���?}���1]U��g�RG�kjι��o�PŜ�x�x��q�����/����o�Q�k����ץ��+�XGcd�����8�;�����ط��K������Sw����4���d�eq��#��Z{
�gLɷ,�j�E�?���̪�H",�w[��a���h���������L<���U���������N�5*��~�!NH�G����L�����M�O:N��1��l�떒G�~��5a����3d!�{;��"��e��sKIK��X����eLez&2�����[�B��ٚ�V;S�8C�l�r}����9D���w}�7v�<����t�f�l(�mMʉ=�����=3�c�'��&�x߈+��IOsi��rR�ֹ�_6`�q����ӎ|U-�^�9`��P�s���`�2~g���>�|�����9��XO��J#��rK���E܉?��SZ�e���/ð"�V�������)q����1��*y�l���-��8�q��,1{r�C�u<	g��Hr/�^����+W���C��:+�nד��gT��dAz�$b�	��^��ϲL��g����:��ރ#>!�`��ș�Lب�8���W�x�0�P��N__��p� %��54�k���s�܉�uկ'�]n�4	��~�&�Ԗ�':-�nw��~h�Θ�@#����]��������p%̪�X�^�����_����D��:�e���u�+d�k����h"g{� ���.�D f��������|b��[2݁yry ����YG�y��d2�}n+�{HdS��#M1��V������G�n�0�T�2<%��Q��y����<���1k���cń�ă��aD��:��
�cu�����J�kv��@�,pʝk�]���|�O���J��:�}!�%i�gn����,�H��s�b�b	E;�B����.sEh ����C��0�]a�<a��%�.,�̋�a���f�K��v��C�?�B3%�_�`
�c5�.���G@��U;���_�+,����`��(�%�z�/t�W��,�D�;ֵ� 5&�ŒA@�p�kL�5�՞3T�6m0��RZ�k������w��,�fNZ�h�G�# U�W+t���v��2�+�T�s�,dyS&�߲I'[X�}�=z}܎y e�6m�G�������n�^h0X�p!��و���U��h���5�`SWh�N*�B��t�-ϸ�%I��.����72�<A��:��vYY�H���Mς��1��D����Jr%�}{w�Е W8�Q�W$�P��(�M�
��ˀ���gOB���?�����^Q��`^��/��}�E�����y��)���{U��ߨ�~n&k�H%D�&gl�aqj�I�%vkr�����|,$�<�<f�,i�:�*�����>���IU�!�jE�Y~���}�L��q�Q��pweM*��O�mG�OR��,���#�^K� y'��P�����?�sݹ�tƩ]����/}��"�m����KK���[�<lQ�xd�	(���~�$7���*��ۅ�_�;�2c�o=��B^�:�d���C(��Q��$�$��^�0�eI�J?fh�\{�_C�؀�Y�(���A:�³s����b9cB�H�B@�������@mʒ�(���<���Kɨ������b�3�
Re;��@�`@@�&�%"��c���������H��^S�V�|A�7̲RN��ڝ�>��AK�D�.�*��<�l`�|F!_Z��&op���I�۝(�	�Ǫ98��fRM��U�1W-K�X�s��{�H�'{��G.ŵ����9<6a�L�k�͜4Q�b�X�M����3����t
kƃ�p��v��xl52rl:R�C�ە����`���d���I�����z�nǆ
G�|��(�i�K��ڪ����I��`���^��{���M[��WuD��0'�~48~�  ���N�"�����ɶsm�����g�����<���	��W.*.�r涇��RMv:I\z��ր�Ir�-��v�LV��d��������Ǝ8�f�^��[C���d�(nC�W��@μn#��ۣ��&�����/�O8?��V��޻qdN}�z?8��`��`g�x��hTZ���5y�t@���
�Ky0j��?�:��6�!.��+rK�u;���y�̼K���n���uK�R�-�jrq�{U?CE�C%�����|��m=��l����S��G�i9|��
����I�����(^��Os� a0�M�g�.9K�G2g�@o`5�>-~>���ϵ�$Vkm�w���<>B�z� fT���N�іa���B�b+2���->���`� ۅo�p?t��>�1Y�%k_��_����L�=T�7����CO� ����;/mׅ�cn��st)F��3]G��w�N��A^�����&�ۙ{�����H7�-H�3Td"��S��$���͉����kMX��v`W�~ �Ju�K��zc���G��;W\M@Kpbo~��<�����l�uع�Ǳ?��A�
���W�C�>�,5��`z$��1��Fn\_{�����p9�]�k
9��+}QFo�򱳤�UC8b��;VWr=��"xR�!���Ǟ�Cy<;Qk���fJ6O��ը�������qdb=�t���$\��H�Z{N��}܃��s������a`�]�LԦ�x�����]�����P�˚{%ƈ+%
-�2����]a�YK�bb��8?"�$�Yk�u���㇐��J�R3��$�d��׿�G�eh�x/������|Ҵ�r�����H�b�͍�ޓ�]�������t"�b2�U1L(�����	,��b��[p��V�z%J�ÿ��n�P�QU'�e�$��7��	a�Q$?+�F�m���|�+�}ה�¡8��%�1g&�+�����*3�mr��y���G���UuF"�N���ձܒ:)jl7%h8э0}�~����#ak�h�њ�߈��@ekw�R�E��g�:/��CFUO�������"��bm�����׉�5��`��ς�}�S��8�q�׆
?h5'`x��i4;6�>spk������ ؉�6"��E1�:4�W����u��2.-��(�~��lj^HRR�l����� ��$[��P��)���c	�h�b?�	i�ek����t��R^5��\��(�4'��)h��gE�Z>���F؛K�m�X))&qI���������W���P��+d~�e��#A݃bSÞ`TPI��{L��+��;ϟ���[h&�&��h��z��%_֛D���F�.��$��S�@�s���Q�V������p�ϔ�8"�Dhl����&��&y�z����V�?�`7R���.�a�-1�RA�$�.@�� I�s��4W�Ҿ�; тC7|����]�/���a���a�E�����~�E )�X�S��܊ӏA�f���S
^/k �J�Z�����+9rd���Z�Ձ���vqv!�]DQ��-�knI��s�Qsu�]�|����� ���vy�@�)��ߝ���R�fl\��j�L��q u�����}�F@����y�j#�I͗Rݪ��J�0%Zjq�cc���3N����b-��Ё=�;�U����w[�S�r��ee����珐�Ą)�:}�����������<�7�]Ukmm<ʰ�Z���È��-m�Y�K�ꤻ��n�́��S�	����kRB��Q�In�����I�����)Z["��C믫H7ʰ,�@���٫~'�ן�����,�p������"�$Y���jÜ�\� ��#�JK�+6��!WLQ����?:
��|o��Ơ2~l�%ÄK~w�_ l�2l.�_ ��V����۳�]�+�} k���*�����-������[��d��%S!�H�+�Ӧ`D�[��+:�e��M-�pD�=I����(��촩k�Bz���)�`w �ԛ�r>q�b� �Ї|��[�~�_�o�4�W�~n�M� �"&�� �[�r�LBA9�ƒ�SYY�ؼ��5����oyB�D��m�D$��%���Q0���ũ���\�D��^R~ݍ����=���m۸��IVv->.�W��O�$���c	x23�&�4�ɫK���5�Z���tK��z�Gr�ͺ���� ���a�� ��(��^�M�Db��Ą8J�G��dY��HC�ș7D���P�Duy
�Q�aR���
yau�����KEߕ���4Wb-��n�]n��5c���J�O�|D�@���X�}���|�(���.G+3��
RVn#`��f��L��/9C�:�x�7V�f8! �*S��f
^d��ӑ�$C� X��.C���3x�ڐ��0�V�j����Q+{�;C%i_c&�2�,�el�B�;�{^�Sd��?��#Ο����<����6�u�W!:V_��^�6o�����9:���6���r������`�~d���shv�ߧ4	8B����h��o!�o��t�-����U��)������X�eh�t�#��	�69�/+m������C���RҦ��ɠ���Ѻ�{�xj�%����k�K�g�xS�ɸcl)T.3.�� %�Ԇ�B�UV�s�����S�Y,dx𦞎�1>>*�Ժ-B�$شxK�� gY�!��I(	(m(i�w.p-�	/�i�.s�9�r��VC&r�k:-���:�Zȏ��9�O�0�6�Do�a�ӆe�~�w����Q�?�RNM�w_ ���}� 6Ւ{�R��g)�)�B9u�,�=��.CI�|IA�a�39�AO���.ՎX�Rf��Op�4]��FpȍӀ_ۃ�����ى)� o[����_B�����VW�V������f^2����SЗ�S��M4%	��=;.��AZL4M��&��2h�$t�:vB���7����QHU9,𢆲1p)�����eF89dj�\���p���]���-]��TUv�ԣ�_e!����~��}����i%0�a���߮c֬�9����g'��)x���zw&�m
~ ��y�;�x.�ˊM����R��?̖:9
�h��B\�1>>�d�2�HB6�L�}Uz4wv��r�iyP_"��ۍX^�8�A�'�a�Q��7�5ߎ_A��u{n �����/U�~�,�k�R���9P�{�U�@��Ⴣ3U��;:�j}兒�騞������#���e`m[����gڗ��] 6$��0:�"����|P5�}s�cT�4��=�q���ٽ��Bn������[t\H��_�Ğ�1��=u������ �l&ɢ�w���v!�����t0k��j[�I�W=��&<؟�����C艼�؄p��F�pҨ��A�
�-�X�Vtmtc�q4���⒀<��)J��� �*�U���ډԉ��8]J�LE��2�f]z��������������"��� >��"�"E#��"]:firpж
Ǟ/�b����/��{�88�nK���3�b1X�@�WY߶	}���C�$���LԂ���ΐJGޤ��ҥ���9����1�Z�bj�>��.)+(�C�ܾU]�B��YӧTuQ��]	Y}�MѨ��Ys�>oX�߅>��3��mz�V ��PB�HDG�*V5��D���&�|�%�G�|;|L����W�Ax�/���Vx�Rvr��P/���o�BՌ��2���S-U�V�����I�o��K��$�ml�	Y��>�EmG��� 6RJ?\M��}R�D�x=�Z�h�d��xl���J��#yh�7��~4��K��SD��Pٞ�*���U�:n ������^;��d��4������e�:��v\c�8PZ���_[���z��{| ��H�}�]���-f����4��J��1�U}�Z+����:J��u��,���/���������i���r����|l�kͭ����-VS�����2q�)N^$�fm�����s�NM�P���[�HE�zY��V1|8�%�.{���k�ce)�{"��t���WjK�bU�=Y�@ԴS_��9�oP���9د4�!�R�?#E8&̾i�0ܴ���{ͽ�P�jTdPn�кG�E�!�/��g5����v��L`�>Fb~ö[���铽s9����:z�!���;�b<g#I����;��fg��-�5�R�uY�O���AJA'��æ�q&vVo�@�}]�ٺCj�<��_(�t�N�����Y:}�����[Uek��J+��Y��e�����^_0��4�i
"z���v)6T�y���""�`�t�՚2$uʲ͑Bp�:Vuğ�O�M��<���*�=@�
�%�: i��\K/R�'�
9��Ewo����kC��t��eH���ʢ�:���CՌ�m��By����g�M.��9�P�#��82�xaԴ=�}y��^V���~Gz-�|Jo�_�3z�� �H��y �Ζ����"��2�T$$h�1��ᆫ;#n�)��P.k@��3����n)<;h4�Z�d���>򐷢����x��7�<�hn8����(�*��J�\�'6$�4�>�3�.��Y���T)������M���S{���i'x�B0io� ����v�T|��hM[Y '��UN�f[{���"Y���V�S��h��  �mK��� k=��(;g���}��z��q��j��y6�G�fNE��,�k��)�52�.�`)��rn�2�=QfD^� ��.c(�� #���x�}���8;��I����H�Q�MS�K�@d4z5�	r4L7�m|�_�K�^Ȭ6�c�BW2w�K�^�����rC�Ovw�a�v��E=�0S��u}�U�R0�M���_#F�H���2�[@J�xKA���z^G<	�i���c��/Ch!�p1%��7V�Ƒ��6�]�����<w��v�+ yc��hAޖ�M���il�@o-"kr�<UK������OD��;��w<��]r&�I�G���2�桖w2ƍ�>7%k�~�q�]�Q����~AhEK�� y��^$C���{Md��Q�G����0�ĉ��7�<�zmNsWj�->>~�O�
q?6>::�,^v�҆��a�+��`�l��Ƃ�K���$�[���IpwHpw�k�5����?sgw_�|u��TG��z��$}����f��w���[u�T�����������=����p��H��S_i.IE����q>�e������g�#��o50�^�t8��l�Ź�mFuH�:�>B�� h3K#n�0���Y�݆կ�ynf��I�Wc��6:s[�#��QL��Q�8���'M�z��8+�����h:��b	���N�俗/s������	����_чX��F$�a�3X�hy&9��������`�r�Ҏ�+h(�g�d����G�@��1�ݲ�;�|�c�l�g�E����E�1*�T�B=̒�ᧃ�IXQ���>V�y�I3�����Dq`�����J�>}�>z�|l�o^�
�7ؚ�g��z�pZ���e0R<���(�����AN.�|��|����̒��J(ǳ!HN"�|({���e����5a����V�C�_+��"�⇔7�[�����2��*mL��7�i�^����"9T��-&`Y(1A?�?�"ԫ��1f���X�	�lT�l�ҹ��:����k�����9�0�?��Ij
��!F��0�N�� ���!/�N���䛦�f̞�߱�\��x�ey���&op�g�!�	�d���[�ؕ�� l����b��Һ>�X�(S.�
�w������|��*��� pT���"�{&E|���`
���%���`L3�Fu~E:���=-��qEEK?Ce�kDɷuX��lS��[��D_��c�g�cI�|��"�VZ%�a�����>��Z�i-ja�}ֽA��fu]?y�˴��r���eJ�-�m�Н��Z�C58Ec��ն�*kn��ka"���BWv�c����:��y]��3�E,J��ͷ��~o�T	��ۨKf�n4V&�q���kS��#U�n@��֫���U�<���8�j5�Y���t���*��6��X#��T_����5����,ߔ%F`}:�d�?�.!C��;����G
+n �G��T("�x�Ȏ�Sy��f�����o���Ⱦ|_vſ�_���K�wm��݀�uc#>�p�~��<|j���Sg����B����>�0��&�������#�OSlB����$-ny��YG0Lobu?�뮡��%Zɬ� &�?�(��p&MڴK~�����\5�:g� -�;�X��p$��+R�sGE����ļ|��t�9x?[H!K��eO����9<��L���B��:�<&|�SmbѾ?��TK]���)
[�|$s8FP0#R�1J���h�lSt��1e��fp�+	�c9T揗�j�`��&`�	D����w��
����!�,��� �;��U�o��iZ4�Ұ�����~�M�y��k��-��@�Z�l������"�6���}9op �0��I�?T���iR���QΖI>
�$9�Z��RXa§�o��0e��2',Ae��7+��Wk����J�J%�тnÞ`�I��༑�H1ǻ!�i̿X� (�/�zS�/��'4�!6�LvX�B(��xBid�m?8�-�8fY䭎y@����o�������a���f�$����ν�or�c֬\Q�+�)eux�[�H��y�������x�̓+vm� 4����=1��b��D>�:hT>�nw_�C#�B?�-X�&�.�=f ��q�����-�2�+�m�KY�H]C���V<���*�ؾ�H�(130��<�W�h���ש�JU��2���<��l5��[Ϲ��'��]���a�zO^�
��(����Ν�����x�d,l�$G�GD����YpݹEa���e��P�i5�S֐Y�^\¯YF_4X͕#!4g'�H��з���R�Ä#!!����se��C<�z}ɀ�ı���3��)Actyy�Ѻl����u[���$]8V��!%?�l,��C%?��k�?O�l�n�B;p*�fl�������BSN<����'�̆����ʬ�g(=��qhpQ�|�ɾ�MRP��A\���$R`l3�b[�ZL[7�?t����¯�.R��
�S��� T��-?�x�$��G5>�Iᡉ`1����:U�,͡���`��r��?ʭTSт�`y6�)֝���1���u\`1UoX-Z��g�}��QT���)���Ӄ����x�i#Sa@�Ai̐R��_)�e3^���T팴��%Lj<�r��4�FХCz�a=0���I�7H��f���s�!i>�~(��n�x��`�?]�0�2�7O_��%� q�a�	^�faK�)���Jj�2��+ވ�x��_��$"�{2�;�WuP9�[��+Gt���ή�VJ��K�̮)Q_���
H.k@�EG2�Y���GN�ҿ������m�>�j'AD}
�E1�\j4��`�]�h�7����Em�N���
���D	��� ���۸2�����開T֏��L�ڛ��Y���TL���2/�'P�_���E��I��Iʘ�땋�z�Hk�I�#N�&B�H�IN�p��̎X�ÿ��m."`��9޶Ԩ�fK�}����ւ�����^�-�����9��%��Dr=���&rRΛ��ƪC��ec��1�`���OQ�2�c��ʘ.�"�Dd� ��=�g��ӄ.�H�rp�5�툆<W �b��e�����"����2;~����:�ET�<�.%}�#EQC�-�+����˛i����f����f����`p����W�w�}�^��!n�)ԗL�d>�A�fd8d�ݚ���B�˕��ڀ-*>��v����+���J�d�����ɏ���v�?m�[���LhB�cgRo��-~?��>+?" �jNtL,��^_�ϧ��8�F�:�hQ[�^79As��
�s*�����Y���d�q��.�ȿ3iL�l5�]�ڣ�WD�di�e��[B�9N;�Gȹ�Rbמ�g�� � %�\��;��uY���̵�2�EY}�μW!��k�+Y0Vy@���`?
�lݏ��u��X�� �ּ����-=��*�m�����%-!��m0�b$�� �8R��f�?
�&>�9�Žb��"�<�1�*�����7�9���:�����+��#"�u/��j�|6ȥ)(�'�<� ;�+7�8�p����~;��$FV)�"�
.7��V�h|M�ԗU���qdk��3ߖH18!�6��%�=�T_�Y��v>���ϔJ�m��`5[���L�,+���ֿ��}5��`<�?�0��0�FQ3~��H�Ɣ�AR�fP���(���6M]f�C\���#��ZF��E.�P<l�J*���S�'�P�!�Q �F�A��� ����,.�klbݫY��*t@0�f�����h2��`&�b3(}����^w)��jx�:�SG����uY8�aco<����S:e
��0����ł7p�5k�"��oj���?���8m�p���	��c�|��C}a5t���S�wy�l��� t7�����r�p�7�Y�v�T7�����D�IG��������r����u�����9w���owfL����=��U��A��s�A�%���m�8�����,��ANJ���|k���Q�("IIX$l���'@�!����i`��N�ھ+՟p�y%\t��ϲ9�x�J/�n�y�Y���J���k?D�Nc헭����hc�v6�c(�ϒ��[{"�[�׎hխi١2=��b&-�ݐJ�$���v��bG\N���)�֜-`9���-�սֳ��HS���ܠm��Jy�F�2m�������n5q%R�_�?��O:@>���h<����ޟ���p�2Do��eV�8m��hպE��ˈ�dn���o���N(0}��b�����YQg	@䠿70��i�]rm@��B8�o]�l��߶���A(�!:?�e���ܙ>��B��~�g2�=�o�����qS�4ws�ig#������\��/x1C'��d��7�[��������U:9�	���G���,�
ѵκ��c����^�L����=�A7E������A��k�2�9(�m�S�4���@�?�����n�^�y��+̡<�+y�;�����-���)�h�n7���V���4��?1:���r:�1)|1y*|Ѯ�%�f��� �F�T��:��eiMLbz�Teꃖ�}����í*�O2YN�ʓ��w�B�K�j��8���.��J0ፉ�P��?*r+�x�9������(-6/��e�SD8�+����t?�yJF�/Z�諻c��k�������y�<̀�&��|>�9A���4n�����#�����
/�ZB2ig+v*E<��_�$S°������� y�FIh!�~�c;���N�b9m&R]W�����?|�ג��s�SK��o�XenOF�r�if����d���QR�����q�W�����g�9��zy���%�ikh�88�D&"f�t�@u!UQ���\b�N�~1�!*p����c�����wO,`�g�����9�)����ʈ2�+�pKp}J��/����@�G�p�v�����@8X>�x⍛�V����<Ux��/>��}���Ax�:0��yR��ş�а՝J�ʿ!�~~�Z4r�
x8�l��h�g�i��<�2	��!r[މ����T+=�7��w&�����Q�3֫�g䖵�|}�^�[��r����z)��pr� 9� ���J�<�����V�-�y!��=ھd\�h��&�EA���T���l�-�8q�M���ϯ Y�n"�)��ݮ�[� T��~�߮c�~;#�d��+�"%�X���'��3�6m-�c 3�����u�j��
:��O���)�`�L�yI7I�U���g&���F��ݥ>�7$�Q���g�5N�y$����q�H�����;������1�Wz����a6�v`3rQ^�(}v4)~i�f��[���_4�"k�Mv��B����\k/,��@�n]���$�%��?�=�y�ϩ�s\`4�h�VSJ3�N�ķ�n�~�t�7�v�]qPD���[�>��Db<�c|H?��b����)A�
.�l�A�&��Ty/qI6���eN�G��oԘ��-������@�l����l��#ʮ�/sa�����2�G@SSb.X��6�ֲ���72R�&�M|8�?�gR����L�L��;��`�L�ލ9�vN40�A��>¶!�������5��K��Ǯ~Br{��vGk��)v���H9�X+��λj��G��ͺ��ȠO����T9^S��i����{@#�{j�o�>J8+_����5>��*�(�y�du����gQ%�ob������U0M�I��!�p���v
�e:R��|�H�I`�#�7��}����t���z�ŋ쀞"�yAÄ��Y�J����3�Q=�l6%_΄7%�mPEE��{�ǋ$�Nh� ��p���(�"%pv�v�*%)�NX�U�?�G ��%�Ҽ���At��P~�I��L_̋��|k��NEZa���%�KC��p*�+�h�|-�'�c�{@�ȵ{d5��m'�����鋀��8�w��e7����  �e��иQJ��+63�H��h �9��`GU9ƒNbg!a���&奨$���K��S#��OR���)�W��u�%:H�NQڊ�K�([�����\��F���������ћn��C�\#G��֒}RD��ZW����Wi�ԓ�f�3z2�*tR#kt��G��u#����F��bM����+J��m,���D�IY4�>�.��'���hN�1��X5ˆV�d�Z���J@'b*X�8��K��9�#��⏳I�^��:)�
��,��_�6��lY�ߵcP*��N�V�wj$��Y�����O���I�!�����}.�c�(r� �Z�j�D;e�D|'Vq8��BT���/�	v� �o���G��O<;6�aU��~�S���:�G[D�Dc�z�D�D�s<&��0Q_������İ?#�Oh�l���7H�JsY��S��YΔ3�.���kD9pYۺ��܌b�8+EZ��ԡ��9%e�ꙗ|�q�Yd%�#��,'�V��Ø��:�V�"�x!|*�	"��k�%�by9b�7 F�2�ā_�'�:=x��S�r�����|�1JxC�p�[�X
��+o�A�2Q������|�U�Ej�yE���$��Լ���%�xF��Z�d�_8Q0���_{�� K��[����S��A���D�����,��2ߥ�?���<#����"���we�U.�_�G��3�|C��c�c�^k�X��N~��uh���aC�m� Ϻ�^J�>�%��擢ּ���1*߿#~�/ϧ#��d3��Ny�~� ��D"�yEO.���U?*�y��4q�ۜ/GU~>���mR�����F�:QW�=aҬ4�3(&L���'�ೠ�;j��ec���LJ��DpAJ���(�GiFa";ƃM�b�>k�����ǠF7�#���θW�9-_�m8��2���h`�G�%������;>���;���'���,�����FZ�B~�A�M�P}�l�hV0��%��:���&�E���+���V��Udq�p���)���iL���ה�2��a�8J~(��Q���Q��jb?2Z�>�T|�ܬ�ʭ�K�`g(1��Y(�O!i����������A���/~xl��}qsm �"|&l��&�+�S�e=~��<ZVp={�����
�ˊO�6�v{�m�f�
>	�CZ�D)u�|�I���u�[����U��*�����6�u�P�b�Y�qyjQ�!WJKr���T�:]WL�P�b�u*��0��ԏP|�B���V���5l��CQG���M#En8\�K�<���r[s`]}�-��Tf埊��x����#+LI��v��v������f4����ݏ~_�TG�kmW
��ǹ�#\X��!UvQ]�Hh�}A�}}�a�,u��ߴ�J�t��X2�[1��Gg�'�(�+��O�^c��0���E���\m�8�/���j�� 	�gvZS��eȺG-���~�Wv� {o-(-
�iq�d�eo$e��WT)UH��Q\�~&��
_��b��
�c:�dq��4	�X
�[��ШY�GU�DL9F�7c?@�H��:0Z��e�`���+;Qo}�O���Z�̜!��/�ܷ�*�r����iK)pB���@Y��2K@��.v���ȩ���t��Q��z���Q4���'����q���M���k�>��ѯ�-�z�z�!�ON=����G�j�!	�,i���;�1��J�Ό���@=(d�H��0�#?�C�Q���
@��9L�|qx �@���Ujc�0�V����c��p�����0���3�A��b#���2ѓ	C��'�T���o���j���(A5�߇�i��D z*c�Y(SN���7�4��v}��6i��?��P�}۩6�V-cK����/���cS��}s��,�P��s:�c���P
��p���)O��5�OE/L*_�h\^��8�*�����"�GG�nk,�"����uxB�+G@����ڛn�Z�Y�oF�E#Vb7jY%`�f��glv�z�?m*c��>��{�����y?�X>#�E�tD���%�� �,X\	��)������|����s}���5��L��hn��������.r�Щ�Fi�%�]��
�9��)���{�����7{<|V���/��S�X3�Z����xP\�����LF�x|�/�h��v�r��q�wV��� �|C�
-<-J���H[CZ��
AjQ[HsH�ia9@-��M?�:Ӣ��8t�]��NE�Ю��-:�Rn�k��B������D�� _b��r��U���{�ٖ�?��VG
l��V�t ���ĭ �-����͹���=޾�Ҿ)� s8Q��L��o��}��1Gp���}�gp�b!K�8jƑg��us�^;����{$^��:��/B��A�(��qy���UY|S=ۼEᣳ��*���f�\�ٮx<��*2�)��#�!�V���v,���bLU�����li��V��Ō#q��
e��T��{S� ��&/x�1O������	%����}4�])���v�����гr��U����3��׃ԋ�7����$a�Ol;������p��o�׮Vz�G��!i��j��z�CQm�>��w~�]F�}�%��(���["� �c
����h�N����0n;�����GJ�=����`�B���C�;NGGG�i�ʲ�x�E��Fj�o-Ĩ�R�=b]����������>��o���g�|0:�o��L�x�z��F<��48�\������x�o�e���`r����rn}�������g�m,���D樝4߄Ɗ_��.��u$�//�b�;�5�O8zXBG��_�8Z_x�n��=.?dN���;U�Ê=��Z8Z�X�	�1O	8vݢ�>?��NӴ^��n�d�;�=�>�~��Y���H(!!��ѝ�q�	1��Zݰ(yM����{��z�ڹ*�@�<� ՞�.��`Bbbb���x*�ӝ�`K��p�z�`��T�E�����;i`��t���W�2#$jᯧ�}�CI�B��GD����O��**p�k�U2d���!�A�r��/���q'$��o��OBQ�4�X:=U�~��,O�>g t3��d��Е���OZa�@SS<ɿM#���o5'��	��%1�%�a�d�g���:p�hB������7�l>��d�W}6�7�@0�K�&�Z�m�K�Ei�
�K���_| 4C��̼�(�E��D�;��[���7h/�BW�6�G���]{�fîV(�-��?���B)uh����`�T��s��u�?hO�:I��:�e4�&9��8o0b���V�\�
)��7U��ƈ�hXa�����%Ņq�> ��
qa����&ؒ}�����q������a��]O�z���?��ɍ�����9���1��Bu���\����#�y�����6�۱L�;4����ٍ69X�F"��L�u�G�����n�~��ܜQ��1��uj�F��G��!��?n`"�O�C���8>))y���=�|�ǯ�ՠ��"���������J�[w��?�|��ZFoYK��)�m�s�K�Ϣ{�b�e�)�^���D���ѫ�V��� |׌l}���$E�NU�תR��чJ��'���.,ņ~]G_�qyͮ���O=0w��q�ވ2����_2qedqB���"���h�2���Q���p�(�&�:��\_��T��d����p�q^�̩I;�ڨ�l�}�Ug�'Y��~�U�ؒ{���Ӵ��T���J,8#�c����T#��h?s����[/VI�����{f�֕s"��sc���k�3P�9��)A���b`����^��j���\�e��6)�n�X5����2y����ҕp�Gb���~-��)�<���}�'rh�qH\�!M�ҿ�D<�;�p����ކ�*i����ŏL*�}��Z��z� 1����9��O/�#!T�Q䁘�%�ci��]H��D�5؋���//Hmϲ|f�ٵ#���_��)F S�1��7�������|���r���^ �ft�g�HM~�>5�z�6��#|�5ñ�J�OMN7܍��;(��ZA�C�O�J� k������.�y�	�ڽ���#h�(���_���ezN�L�+���G[�8����z-�ڴ����~B��N��O➧�i����?&�d$���&�U
#h{���o�}4w[�Cƍ�s�'�8�ˀ/٣{��y�r���怵@�������S ��*_������N1"Lvk=Q����%����hP!po��aBy
�x�Ƽx{�ݒ~X!O��!�H����卑ýF��$���iM����j6M:1�-MP���c�Ԋ����av�f�iD5�@����t��f颪�N�x&a��
�u3 5~���rE���c]�ky�iF�(�S��ї�\�U���>j	�;�;���0#ٌ��T�8ղ��Ġ�?!�o_��u��&Y{����%k��\͖�'F/'�^���&�Wl��z]�t���(�d7�r��vY��0v�@`���lɊ*^�����圍�\�`����*�Ql��l�o�\Ɂ|B����̕��YZ���l��PO�XI�s���d+�E˙v���3���+f��K5���o	�g0H�^ �-�Lu.]�*\�������Y�惍�r@cBH��́�pL�d�e[��:�]F�����V�5�W��C]���p�E2�шC���Fn��������C��]GD�ڄ�����M�b#y5y$lz����e�|k����kۑ�i�ʁ���.:��P-a�@$��R����u�_[͏`�1b:��@nK���X)��a�M,28��[����b�/��Rﯶ_��Yh�Xǵ��:�}mt��R��m�d�辕H��d�d&�lQ�ϡ�<�*}�
��VE�c�E�Y��f�	�-�M�旉b��*eOr�?me���mjڪ�M�����7㨰�xnd/�i!���g��a�N�E�p�i��	�#�p�,D�H4���ԦN�X֎$�B��*]����h����=������\��JU�p���c,w�vz�
'�����)�$�~���P���f�4�v�b�S�E8�F��k�����y.��D�r�;y�;'*��vr��:L�c)����Y���0��A�]N�O���l�7�|Z�]�^�J�|�^��u0#��o�]�bF��psP�4�����^�-�Y��,W�/�0�� ^��CbDX�J]n�dG}u�ޣ?�@�l|gh�	���ަW���ws�������Sh��0�㮍�4a��uH'E��
KM��=o��������
8�JV�w�+M�
?����Bo�/�`<_l)(χmV�����u�aa�J����>���K2�A����s�Ʋ���hT��[4��5��F�&̆,����_"Ｚl��ȻOEMkx��M��	v��ϋ�	���y�����Ue�L�/ު̋�k�-JeA��W,�~�]a�ʚ�aCI��%Ӎ)%�����V����qM�\�2�*�K�rm��h���pfY��n�x�g�Lڮ���_���*./7X:@����0=�II \�Pp��Go��U���B�_�&�Y�^��b���0'o��<02��*-I4%o���{_�~�l����y?U�V{��l�:6����!�^�kߪ,�q����V�[��V%Dć�ٹ}�C�v�l�� �b ~�l�ݒm}ˏ#P����F�S�{\��;0-w���

��n qZ�kqr
��t}+4�v$��I[�伕"���
��KZ����U��$�+M��D��c��İP���֗3�	���qZoGX[�ig�KO�++B��h �B�����f!'<�>��#� \1�b}�SE�a	���&eq����~���:�JI�&���ldNd��	��e_ݦ�R��J��<�+�����w�����$z�{-�ܟZ�nes������E�g��jT#����w�wN$,��;?��s�%��xFh綇Jw��B�Q�4g��ʙ�J�0~,0�\F�X�8�F���s���~��&Ɉ�6���:���g��.qEY��H/�~ɽ��_��B�8[�nR2�}T��lـ/�o�"="�`�9�����ܲC���)U���d��\ѷe��i�IT.�ϜR,Rn������=��D�)N�Dh���Rņ�0Z�X�����Tc� a�iЊ�	WQa1U"kH�;ϧ�/8p."�F/���h`:�r��H����H��#��c3�����ϗd�>H���c�>Q�:Q�B�Q�_`���=���<<@�r��Y�q�~j��au>X�9��1���~��]���pS7{4Yp�zY<�z�ǃ�n���o�	+%!�(�H7B2TSFB��1���A�_�v��(�]�p���`��z8~$F��I:��Gӂ�:�O�R�B�1��Ge�3qrT�b- II}L�:�T0�{gD�R���`�%�g�^<�@��5���p��㟯���p�r9J�+~�`w�f��8]m��S{ �'�����n���p�����a���ͣ��R�5����� F���P��O#�}}/�9k4]ҮK
,�Q$%}�/�����c"�׳�p�3�����qS�ǋ�1��N��q�PN҈хm�&�u�֚Dp���3�*��l�-;�-�yԴ�4�`aYo�����6��p���sJE�gMr���?���5˵�@�hH�/FK��ٹ`:�\F�����B*�F9.Xݼ{RQ�t�|Iݙ-l2J�N�W!]��;,��̡�Hu�C��Ԉ,{��ft�g=������c��x��^�\���j{K��6�0�u�Osm,F��nO�:C����_F��uq����:XӪ��*33R���g���
E��	���;p��a�qcvښ�n~M���;\��~-���0<o���^�g������¹���C��������!�Q��E7�����aΖ���6��`��ʺ�˥�G6X��̣��0{�>cT��B>5��4
�%cۖ���=��C�;�o޴M�_E��c����RΖ0���#���>����/������u'i���^a3(I]RETb+z�ʋGԸM[�#�Xഝo!�Τ~J�#�r�$��|W�Y�43D�c@t1���W3?T:m��R���J�;Բ����w�`_�3�%E�{��a{����%�z������^`@@j=��m�q����6�g�B��k�d�	����=ȁ��4�͝��i%�j\g�����y��U�$1����jqs�Y'�=��m����H�I�����{�ٟg�|�]W����;�F�g��� ��z�5��NF�UC�t��2	�e\�k���i��y�	���Ӗ3׸o��v��/�SHS��^m�m��G`�61�.ҡS#��M���|���c¹�{!�������1��A���I1t���Q��}���_��@�@���jG�:��yL4ҷq�#�xVu��t�[h��4���m�l��&,�_V�Ǎp��?�f�0A��(E�&u,wN��:=oy�{̰nd|��%�b�o �UB�:�����]�z�o>��`$���z������j�k{E=Ů�CʂI[,���bl��ŵ٪���՘�锨ܑz��*�6���ՠv��D��̲ �A�
6��`��7ſ�Z-���R���fݘи\+��#�;W��(-X7�C#>	��5�B�,:�Y������n@6Td��o����c��:�}teϜ\�-��U��������v�Fk�*������I�1D�X��a�E��8�C|W;Q�#?�TkB�TEF(��+ʔ�t���XO��j��[H�^�0L�\�`�me+�|{�0�?���c�PdzӀ8����Ӣ��pp^+�S ��e�Z  Q�R9��{\�	��n�4��/K=��`t
�MJ}=m�J�� {z*�4:ΐU�lh��/vL�i����{�UFO��n���n����j����%�b���2h���S����H~p0'����A'�y&��������p}��<l��z2�w1q�U����m�k���l8F���ՠ�F3D}8���v=��]~�xq3���]~��k����^���Ъ�U���
�r�6���u.�{�ڧǦ�m����q�Q	�$��R����N���[XLC�7�ߤE�پ棢��D#5����4�#u��V�x��)ҧ���]��[����XF]�VC��;�o�'��a�*�������=oVf�<_���\׆���0�8�К&�� �K1�����5�}�OS�q���[ض�)��xhD�{eff��;��8���Ь�E𿛱,h3w_bΘk��H��� �48L`�>}6�#�,+�(��6��ʅ�vB�H�3v�Do@���T�x�jv<EP�iS�^}|h��N�Hh����G�
v�Y2���
��Cz�9�_���V�vI({�v��`�2��Y��K� ���}}Ԋҹ<wձ�{s����RsF#L���@,���<�B�����@�=��#�L�"��`��2��3N�La%\��� �d�:�VӋQ��6!�G!�mm��f'Ċ�GT�+U�ܼ�HX��ñ��Ϻ
*�B8ۥ툒<X��Zv�h(���5���x)u�a�6�����H�����i�-ue((��ܲ`rb�q���`��L�����l���U�_B��Ea]AQ?������XʱU�}���0�Va��a����]�e5��u��D>��>���e�g'�?-*z�?m�O�2���D`(���7���M�!j�*���: _�T�ʮI2C�K����\kh�kWD�Iq�(��`t}DO4
�4a6��;vE���8��H�\�H<�C��B�7�N���,7L"��+*��k�U	?����#�r��R��%	��L�k�^oЗ�I��A.���=7q+�@5���?!z�����~o�M����{�EL���W�-a����E87C�=Q�S
$$v��]��fE��̔�֛��3=B�����Y���p��: ��ЉC�'����2�Ь���8��Q�z3+�ذ���zI`B
�y�P�kӽ��xm�Ѩv�4�QOU�[�9�3���1_+����
��Xz?.�!�$ ����<���5���������
�|�DCۙdn�Cd����582J��sq��'�ܘHI��&V4L)�:^�l|V����_�S���$zg\7���?�B���35�,�����B�Ӂ[�,/F��v,u�)�p��q��S�pe��m��q����t7��"]76��g�QE{�X	ҩ	`���:NM�" $"{�b_/�bfV���I��:�KHۨ/�����iy��vI~d��*#p��Ō��П��$]�ݤ����Ӊ���<�w�����p0;.�qI4�^a/?��K��}���j(�&'&�L�7!��SW��4ˡ���2LO�%�u��sZa������P�z����Z�ä.��Y�]M��4[CE���i�L���'��_���<�.7g���Ht����
т������,��o26�h���T�Pix�0#>��}j�%�	�F��!���Ϙp�`D���=u5��hg <O/.f�_X>�~?����d�U��*�\8��0<�rs � "q����k�?utX�,� ގ��-�����r��A�Μ��`#��QÞ��O/g<���������-�S�3��A���ߒ3�`Ng��e��C'���te��P�T�7�/+�����k:2�D��x�IA@<o��'�G�H��"~�&c^���]A��r�L���iM:���7�'�`>T�m!9����X��������������Ȟ�΢��m�g���%�]R){�@�>����˹3���8�>E�<�N��þ�����L����X�U�~�y�ͬe!��Se���XF�}ɮ�pF@J��ٯI�M��BQ�@�T�
��ΐ&��uO�[̲�J�2��(�����Q�l����jAV2��%&]"u�N��ؚyr�qa1\��X���#�AZ�b�Y�$>�X��LH��dn�e�#�&挀#ɂѸ3�K{�K�u�9K�
��---oh�4���7?�l�� �,.-,�=%T�t���z�%~���������{L$�Ղdɱ�B
�P��j��
�׫��$|YǕ�[q$W�ĩ%
B-���КG0�~� Ksr�(w�y��w.S�-=���7��u*�X��m����-`X����[��k9:��Mw����Pd�G��$'���3d-�L�q:QYO��i~���Հ�"��E3mAv	�P������3>��5��[�����6��&�+��<�9���p ]�7+��l�IeŜ��o` ���� s� !�p�"2&Y�UV��2��P�ٝ[�X���X��!"HQ)qC.D2�����wB�.U��~����� �h :���@��M�x`�_ :�P��%�M��*���!hנ�#�������Nb���=��+R����T[P��4s.�$s�Q��ps.0�$$˷g4��ua�~�Z1r!���߭-��dPw�v��F`��p�`~�zF��/C���	˨Dd��t���p'��:&���֑��ޫ�����%��5�.��N���"Y��#�,���rl�8=Fy�Ъ��VoI�P�q��1q��9i��x�*c�:�?}.���i8����TAZ�D`�V?3� �Ve��&����T�G��i�lKk5w�O��;>�$�g6F�E�3��<}!V!������8����l]C!�p�����/4��w	�,@ᮅN� �;����޽/��s>�+c�n���84�A:
K���J.@y脻�o�{��L' ^~}�P��1OK���Ru���<#6?�z��e��c_Ő~"`�YNɯ�%�r�62j~/�Y�ޭ�+z������O���m�Lx��ٯ�A�B�6�+N��ڀ�����#B�e�)�]��ǯ�8p���˴5�֑r��{�<��?`�"�V��_���ݭ�k�$ǘV��{����z��D������X|Ǭ^%����*���ؿ��blJ���Y,�EY�AU7 ���݃�_@�Jl�jTÄ�\����۳ǾhB�u��!�����]#����,#$jƔ4�Ղ��ݪ��wg�pי$��sZ�qp3��g
q��0а��8TG���;��Q�d����1�odmDU��!m���1��T�?���_�Ѳ��%�)����u�����'l�'v� '��#�}��U���ٴ`�5n��<O �En�[�M&�6���c������n������#�*y��I��_`ߥ���f����V|ܠ,����#p\�۞E� f�jc@d�;�n��i1i����LB��<��@Ɣ�5���ؘ�l��
�R�<�uD]�����
�/Q?M�l�����3m���5����e7�E�h+ܦ�����ak�a�|�Wy����������P
^�{�;p�-tFH��A�$����b�4�/3��RX~g�=�T��+�A���O^��w����1h��q͞Ƞ�[�B��_��Jf��&���9C��X�.V;	���Я����i��hl�}vơ�^�����篫ꦯ9�����ϑAX'�X�7
�yr��5���� ��f�@b����ae��f��|X�_����8V(]���y�XT�T`�)-��Hz�3U�RM��f�B1�o��Q�ӡ�*���4��7˥��٣�e��H��@Ѥ��s���y���_�w�:�_A�9�"5��rj�����`�����3�|���΋9���~���_��|J�dҖ����1�B:z����\S�o�XF����A��4�Eyw���"���]J!���3?zg|�wh58���|hDޟ�n��x�9���v��Ʌ�6?���j��.W~�Z��Pq����yU�g^͓�^cX,ʰ ���M��|:���.(d_�qz L��,�<��'�GIkcl�H?*x=�<}�O+瓠Hܑ4�R��ءq�x�v��ҁ��ޗ���=�qG���$���[4*u��T�?M���D>@�՚��	�6����f���������yRM��Pr����9"�aNO� �]��}Lw�?��R�p.]>�z�*��$vΤ�HQ���cJ�2��Þ���\��*ʹ�
&f#|��;úђ���EN�F�󛻸��-`�s^�}w�t� ���;
y��"��)x������":&��Yi�H�e� h�[��2"�'
_��>��	vHɴ��еlO�]b׵pgjx��Q�������	
��p&=�=�g�T�/p�o�X?�b��łB�!r�Y\=���͋=X���[�
�R�y3�b?�l!��?��v�!#ⷊa��7^&N������l3���ʓd�l��O5�M�d&�C%�4����s9/_ݮ���=;�7r���񘑏H:4w���01�j��F��+N/B�����U��y⏪ɼ!�x�r*���3	�AH9dA�j���v��>�;��x���%a�h(�S/�r�_�
�$��)��O\k������ޠ��rXK��9I%��K�x�$�BzʠI����q�`��J�q�$�w�^m�uw�7���A����x	%*�S���L�K/�J��-F����Z$�������Z4ZW�L�}Qtw^b�����QP.���8�����c,Oaw0����<�����]�LyO�<��B�����rKlmUA�C����+����.D ����A��M�!����$�'iz�K����66+���fn��v���
�f?wA���Ԕ&���op��U9���W)�`v���fಶ˯c���>9ro�����J[���-Px�WLAّ/G�����V!vf���֌�`�.H,��!t�[��]�r�^��B+��.l�ޱP��6g�O�à�ՐF6��g������2i`�l�<h)71&5<���Vײ_�L��=án�8�C�6�J�N��47�;c���W��E??��k�Sjɬ�0=���4�L�x\;,yO,Ic�ܯ���;P%��{�|��Ǚ��|38��i�yv| �x�t�L��$N����6)lm]�X�6����sk{>�-t[`�P��[��Uc���zC�j�pq��LC��I����a��;�,��Z,��Mך��8h��<BFq#s��"T��~��.��˞n� �>:B��oN���T*��L�����\�"��:����/���"ą����r���a#�%~�J$lf��Fa��vjȝ--<L�a�60!��y�J�L��h3tw/���SE@7d)C�d�I���%��B��/���[wh0}�ã�l���JH�Z�A�r(�^��g^/����W[��8�S�0����gr�G���Ʉ#�e���Gq2�X��Ш����{��D��
�[ٿ>�Q��pA��m`�������C=5�,�Y��96$B�,��A�Q�v��_߸o�+r�y�XG���p�"�u��3���)��t�f:X�QZVz����_��|Hz��$�C��L[�؅��U)�)e�s� �H�m�n��uA�o�w��B�A��?ZWWy"��*�d����(���G@���+ln�˻��Z�8��M�(>g�r�qr���y�.[߿���]=��ݻ���v߯�׹��֜��6�j��1��$���KTm��3Qܺ�����X���]�ee�����=� �z��`�}Ӄ�x�EN^~�����Z<t�������J��tM;�K��w�nf������,Z����Q*2�F�X�Ŭ��XZ��:��A��kw����B����0�<'��Zk��p*[����3Q�v75L�3m]o5YR��Gjq?�Ő�o�G����!��pD�@+�̱O���\����� ї�p!T��T+U��	�2u��}�%o�~�B��G:�U���O���B�S��߇���33?[�kl�r=;g���؀�g%�$Q��k�&��%��}M�4f��\Bz0�C��_��-������aҬd,�
�$J-M����&N�-�ࡋ�GǪ�9\밤���h�bSHW�p��Q<�+i�1��HE��.Eɣ��J�F0È�XD���*~K����.�KI�p/�s�'��hWg���uw%S�Ǒ?�Щ����#
V4*8im� �ѓ�-Q�6-f4�˸q�T�/KC�=����$q���J�8f4�b8�T� ���V���N����ن�G��$�0D��'�r^��W��^(�VF�����:4|�W8����n��?�ڱf���~��*:��Ճ�N��{��+�8���V�H-	8��������xj��8`V�V�Rw�	�TC�Fq��B������9[�	j&��1��a3��IYf�ƕ
7��]5�e�T��?Q�y��7|�$��Tv<V��"�UB�L�;$��\�r(���`���8=��xx�]��WH\�ӄ9{��u���%��F�ET���kH�èFߞ�㍡w>�o���L�f]�r���EKp.����jFaq��J��
�!�#��������'B-eZ���.֤��c��*���)��� נ_�O�tv�>p���o�f?8b�9N.1��MUJӮ=>�n��#�)
?���ߖ���D�~�a�Ȁ��S�<�J�@�Ջ�k.S�gF7��2��LԷE��[p�������ff�;/{&Ip����!��"v����y�-x�B����h~�4�cO���� #>+�e�gO�ꎿ:��&�M�;nE]�D�xPfI.��pұ��0����#|�Mw���n�>3�N�ڄ�R�|).�H�o�������
��łs"9�[��Η�"u�Y�����~�Ł�
��P�^��e�������rlj�Hf5�y50�X�nV&~T�ǂ��6D���}hP�����"�yՀ����И���2������4WBL_Q��d��*�����{��� �b���[�oE��Kb���/(��j�4)"*c�}`�N#�ia*Sa��B�4>�!K:���u�6#����v���N�
P>+#E8z��1������Ћ�_��IG�[P���"�>�ҋJ�g��T�cAu�S�,u��F˕�!�҅=�֜%W���ɜY����������MxH0궾]Vg���V;ax>Q�	[���c`��nT3-��05��̈)'�g^�����z�/)����6�F�9�[c��X���)�]��4���\_�E�ܩ����Ub�X�k�Q��>m����a���jZ�����kWp\&f>��܏��¯9��̸�M�nuvy�\oaׂ����k6h4�2龜d�j�H��k�,qXY�@
Ƴ1�vļ����W�iR%S�MM/L�:!>y��I؎E�&u�)�T�J��s�ⶌK��F�AZQ�|�Ɂ���E�.fļ.�.?r{de5�י|>�ޤw�џH\*s�RW\���YS��F�7ʤ���ɛ!WbWTX��%�b���tu�.m�Oc������p�<��s��،#+D�>��-ȯ�
�,o����4�]�>�Q�:A���
�K�� �&�XA�x����;'L�,勱�p�!��/Խ�q����/5/g�X��X7�C{h�0ԕ?�I�b@���>fii����|�
���$�
Ll�Ç��� c����bs{�r&��[��`YҐ*�V���q��o��'�c[%�V����g��s�����ś�_��ə��%�\U�%hM�*������A{�xټoc�=��
Ib�)��ޱj��
3i�:#�S�6��i)&˓�r�8)ܬPN���C/�������@�����g�

i�
��J�o���\h��S���0B�j�o��@��%��4��t&i̩dJa����7�Mw�[� �kׅ�ڸ,ʩ�{�ۮ0��41�N�5{�m��ۀ0ۇ��C"���J��:�V˹�C=�4��b�]{'~	ou/(�E������H�3��Æ�+e|�t�
��PWîWf�)9�uT]���bh���k��aK�����v��ωZaʬYB���Z��9����8|�W�O�C<��UA*.�h��ō��7��t�ȇJ�u��>.�Ȅy���n�
oK��88�| ���!��K�G|��`i?g�������<Ǫ��-'"���\V9������f��a_�~^pt��tp[�)�+Y���W��$�9�4�"hV��<���u�W���d?���c���71e��Ep>�'~�y�j?�2t��D4vE�C�o�:4���K�޽����p��©������+��^�B����F�"�5�*c�E�UU`�O�0`���O�nI;;O����<8$CMc)N
]t'�Ė�פ2���Լo�?��S!n����GC�����hp���36M[X��h��M��'�#d�o���IB��M��j�3_e~�$}� ������[�x���=���}�q(sz��	�0���`�G�i4=s����޹c���@������Ԯ[�������꽼�9�)�������g0%J~I)E�dݱ��������#c��_7F�I��%��D85!�z|޴��v(�vg9��>�MЊϜZ�yx�5C�H(Q��a���m�|�	�i6�a�Wu��ڐ/�D���2���g�Z����y����z>HAK�,����Bm���'��Lˑ�\���Ӏ`��^BEPr���r�}�-A��"6j����:j����(Y6����?�o��(6Z�Fd�/�3�^DRZMT��|!>
�(�K?BP�6�u�����o��D�%q�G��+.P#`��uT$i���(�V����v�#��ܘ �"[��*�mJ��� 2�9��A�rp
��}����-�=�E}�&�i���}~�h�m�3�0��h<b�ks�����A?����`�B��"�ԝ!��}���z�@|TN�PH��9�əh�#��#ۼF}�3�v���_i���u�2���ܳOo���WEEE�ǹ����ۓ�V���RPH��P��CM3�%�^?7�oƸ� ���|�:��e��3�&��~w׷�M���/���W�LH$>�嚧�^�|?PZ�ML����O�c�;��4�IE�I�:�Ew�"٠*4u89�`j�������\(���5��%v>5ؤu}�Ghcj^�`N�9_F"ŕa6 E���[�k�N��*s�*��M�WjQ�?B�غ��A��WB����UAIl&T��:�W?c����
�l�;�R��OTO�R��,��1~���^'�{H�Z�&���מ��0oG���|a��3]�㉰�8t�i}�6���Ye��.��%�"��-.�� �0�t�K����,��:�<��^,V�Γ�My$�E�c��:	,��7rWµ�)����4J&�����������`��C䏏n_�;{��<��yb��0�����\�:&�p�SJN;@,�W8?�k�i�Q�c�{ �?�S�"�D_�>��K<4v�%��������f\�b�u�I�d�����.H�F(� k����?�O�T�_��<j);���;W,��vz���m�o����3a��ȷ6d>�~�ME��������$��PV�!�����zۍ5��3�s\Ur_v8$��Ex<���[�Ȃ\��}CZЧ.���Fg��2%X�To�&l0Wx����X ::�N�w�G�c�U�H/�6~�^�HU1|��������m��j��Wᠽ:���.0g���N����`�P��؁�a�׀�C���!b�J���	��p�I���z)1���<��Hc����
<{�ÄD�i	ܜp+`�;��;���?�@�7c����-��R��Ů	ݩ0z�?�9m|����_D-4}"�?�3�D��3f�k�Nh[V����c&���䅉y��v:!�b�K
�"u/U��Y���zE�t_���ܞ8K�ޚ�m7�����t&��3����&]Z�H����wA��%�
 �a6+�\D����\��h}�a�����B@F.[m�=�=X���0�I5���&_R��ң�@���&� ��8��;��+^���
!�XB\�|+���BM�OQ���Ͽ��u/�RAt�Ңa�SÆ?��d�wC�R�ޏ���]���>���������F7�����ƨ�̦�Y�ݲ����t_Жؚ�y@���㋐DI����U�m(;�;a������(�������`���={�R�
g�mg�E���縻�a�ƅ�FÄ�w�K�KϢǺ���kδ� �Z M���%����K�LP��������8xc1��vE�n6��b�����?�<9RW�|�m,CYj�2�$~�����a诪\�qx�Hʲޓ�<����i����M�X�災�7�ct�b;Q�hr�].59��2,��j����4
~�)�s^HN��?/�z��Y4,����_�jC�/���<*���!߉�~��v�ȋf�^��!,w���L� �U~U
���F�m��7؞�� r.+%��"�!�+�`�~�8�F��[��=u�T��t'	�#���~2{�n�Gkg�~����o,@��z�*pk�P��~��Dđ,G�X��Jb�w)��y�"=��L�b>a�,��/K�W��{T%���yQ�8����X���Y�Q�6�Sy-Q�Y�ڻKg�~[s6G��[��dQ��q�=>{�|`�����c�N��N�%�O�qt��P$��ǉ���xh��坹�8�`G����ޚ�M���T�Y�\q���y!�㎑d�\�R?\��Ó��~����a���L�A:���k¿�rK� mc~'!!��.9T�����.��D;ȏ/�O��b�NO+kc�oN��H���/�n,<C����6lSd��[�s89�2�c�'��Tb�dL�����s�~������+��"��"����+���v�3w����+�!�Q�ݨ�d�*߰P-~�͢�o��;��w����^kw�OI��j�B=�BP��iO).�f�)��� A�Hz:�i)�F۟��a|��֙�g��|xM� �_M��F*[�Oő1��Q���2A��~&;M3<W��wj'��V���`��(�~}��$Lͬx�`�0	h�n�2=w�����!n|���P`��ԄU3q��=��D�m�ʁ���(=3��kt��9T"�鮍/��t��N����ì=�f��J�)c�ɏ>
*���f��RV,�E��V�4Sz��&^1����4����֍\o�K�y8mU�i��FVb���0��[��.��h�Ǉ���~2M ?EGs&��ps#���Բ ��S X�`�KD�R=�?}���H���Hx�w�H�',��@�L�N����xB�X��_# !�	�[)N9�G�e��%�R�
�����N�cb��v�VU�>�/�u1U�ǓڟX�͜�7����IPc��B21�ɋp(�&gx�]T�H�������i)�ވ�p@ݩ52�R�n�LLȤE��HZ�9���B�,k{�ME�����r���xH3C���*LGKFդ(60��T�C�e�H���g���$_L{�3�m��1�2L�}��1�c��8�AD�F��b��AU�B&�^$^	/���
��z�;DUR���`d� E��x��f�>�S���z���.��a�0|�����!�<�������ˠ O^Y�@q�*���w�ce��Έ#� %���4�őBA�Z�e���g�IĎ�!lX*XAb���҃؃mDLDt��dU��}�$8>�E�#����l��-�Qh5Xy�����$��2��	}1�;��N���t�6+\����o)��^;F�˧c��H10�G��Bw`]8�A�_|�0��ۖw/ʒ	ߐ펄��:�?ϑD�����`�CTD^hs��z��2,1��J'�thH阺.A:F�L�32��N���ql~h�U���WF�M?#cl����Ge�nS���X_���7(�g�� �9�56��}�F���(Q�o��г�	t�]LJ	A4:�Fi�����4�ĳ<K���K!�ɥRH��R�{B���u;,�
Z"���'I��N4�c�ܮ��-�p-5]#�Ή�4�{�y,|:��I=��Q�A�T���ϞS��%����uU�z�B�qĂ�|��!��ް�A���(cx�4�i��%�jfE�&*m�h��$�h��_'�5�چ���g�v	L�3�n�A�~{L���97��, I$4��Y�£��~��ʊru�BI�yZS.<4���I[�\2�Oɨ6������}�j3��d��g�-���v����� "�m�����aY��o�z����3���c}R�J���=��tö%cFP�{]�Q!Nc�k��?>��=
�	�M�`�n@�Y�敶��L���;�=�J:΁�~�V�N�d�ݪd,cߊ�&�������?���q\�.	�8�n���Ӣ����j�W�w���?od�3�P��j0�xHP�H[����/�6"�R=@`͔%bN�����?i�U	�#w�ئ<��(<�[���"`C_	FimIF���iE���::�l���Q��	sKbb]�%VSр��=�;�ʬ�O�%U��&��/�v "���C�H��j��Eğ�-K�A��6�_-R���9h�߈��>���W�z�|�2|������(��}�G��u�y��8��?��V��f�È�;
��OEMknR��� PV�C*���N���v�|x����楉�_V�W��Q����s�0ef��N��}>Wo��(s�����Չi9� Ż�x6�웢�"������M�L�B��Q��W3�
�p>�_u{i�21Ɏ9��2��&mv �I��_i"���h������Tj��U���E�ș�O��}��fv���{�bd/�u������������d2f�~��������Vs�v�k[�}����,7� �y�yO�����D�K5��%�ba(N��Q��p��Z��_۶�Z�]����kX=��{9�Y�v����nQ�6t&Doq�X&v���Fj;��[{���E��j_Fz��(,?�M�["�5�ԋ��w����j;^x�?,�A��W/[�.�����r�������9
�ǅ�'Eu(������W��R�����
�xdݯ�ا�y�b���q��^i���v/vKZ���X�%f�"H��� ��[Z����Bj� �N]��o��p*5�7�Ͻ��P��뻳���(��U�{YS�0��؛���[��[h�O�9��T�֝dy��۠'�&z��5�^Rsb��5Rqi9n�+ޣ�j+n?6?���0�b�Vn/bB��|g�<��SG�Ë��ͷ���"F�t�;'�]��yt��l*�.�]�֮��Œu�ݩ� j��M�	�(d��ֈD��5��0U�Z�PDX4<'��A�p/L���H�J)�e}_J�	=�����TKDO>Q�.�ь��xп;ڶ,��n�J1�.�3�Trz�v±�B��F��L.��*}�w�����<��3b����e�/��!O�@-k�T��Z����-�����F���J�c��v �TB}+����r5j���c2rx�$vQ�!5^��v�w߮�xCM��vh:=;�+�=ا��=6�ժ�"2�HxmϮ��BO㐹+�+���N����O�?�	���G�*`��"�R����[��;�V�Vcg1�^
�����5�����|��.�Vxi4韥��}J���@���]�o�a|X�}���!�|?����̙���p7���`�3uuH�\`�,�>�ΜҶU�Abo�+�����Ӫ��s�J�I��r�����!W��WP�k��%��2�Yxmf�6��)�;9�^UUD�	�*�a�n�Qr#�{�����MN8K�w�ξ���l`��.�S���8��	��3\����r��2��ꔿ�� �3��hА`祚���Y���6���L�XV"3k)
N��.�V�
��J�z|�\���&���gY�q��aʫ�q�w���p��ŐǇ\C��n�fc�
v���⪦���pI��1FC�.��t�ޣD�d������s�/�c�ҼI}b��r��Ȩ�����k2�����U.[��Q���z +z�/�p�q��c���s����}���u�������l����f�٤��8��"��O{��o�a@f�6���	�����I�^�r��$?k�7��^2���"���ha�R��玧�I"�J��;;��o�����Ӈ�_w�������y�<\�_AIF �!��]C΂�!v:?:~�p��t��PE�Ƙ��o� ��æ�K}������q�Rn�5����ջ&=��
���D�xN�(���~��G�!�"�C�m/1�|~r^�6���Ɏ��tѺ��
��{ϣ=�;r�$̋��[�'��ِ�i�G�p�yN��#9�ҽ��;Q�!,�{l;P6���?S$�B�Έ7��J]qp��{�8Ch`&^���z���&T���ٳ����;�O��:L�8i��%#	�ׇH	$�a3i鲑Mꅓ�)k�t��s����u�- �#��FՌ��-
��.+!���|h�B�
��������9�DF�'QG3�����G��xDP₣�;��:�{Ѧ��纁C���S�6���� �xQ��u�^>+d-x)���e�G��]�{��X��� '��f����݂˫��h��uԼ��$�	O���YVL�ayt|�|��ѹ��Y���\�!���,�$t����]����ć�/1q{�c�������O�t�dj�vA�	�{�
�����8b'�O���#�
�o���*�B�;h�ET'<)K?(�-�_�?s�P��%|���-)���]����X��E���}u')��u"���Lu��g��OG����|�i�`1Q��	m���l�)ꖑ�������
�ӊD,:&�{�H���s2f�#'?kۊ�+g�*���~����Bd�)�%n���`:sI���32�����a?*������d�&�l����T�|q��ߛ05�����Ԙ@�q�gZS��M����?��7�U����9JR���	$Â����↬��Ï40�?�h��@��o���wg��zza�0�5��vN����/_P���Q���
 ��⒨�%��
Z�W[��(�
�;�џ}�2���EY�c�͍��d:S��"e�R<L�e�@[��DdgAf-H��3:�_���a�BCK�EZ��<Q4~�U>H��/>�3.�z&���/L��D�9���-��X��L��:kC��[�$�q���w&K_�s�6?�)���^bP���i��*�'�g�<��HL2}����UF���PIox�c/��\f���T	d�u�����\1�Ov��z`�da�FR�2|�'Z0�"�oR;fn���3�u7�2�A�+���b�kT�՗֐<�\����Y�$ơM������Y0��a�aL[���� Q�����j�5���ؘm|䃡�aX����{�슣VO�ڵR�?l!�1w��{�Z<q.x�,a,�EY�<����+��fP�����Aݝ�9Rh��Y����1�~	�.�^��Rs�'����0���D�q� |������q!.e�oY�_QѤ&�g*�J��������L����d1�>�(����|�up`C�`]�k]*���>��=��q]������޾����vz�Ƽ�H0��Nc�FQ�/���^��ܲ2mmw:J�?��\��!e���ϳ�q6��B�E�g��C�{��,�c�x䦗��2�8��@~Z�@<l�>�d�rg	.^#��<6���ġ\�7�s�0ww��L��|5��)�nq�kD�U@[,�	��9#���dКj��q��ȭF��eeq&��]HϘЁ��`���c(�H���ޡ��	�\��j�͟ɛ�5�F�ުR	¡H&(���@M���e�P�ș�I*Df���ޙ'��7�M�ί���o�給���g�~�Ukѐ�LBz/�kQ07v�:��1nē��U�nA��ymT�4��~�L�"����r�3���R�Q�����k��o��iˣk�H[T�����%���hR��ҭ��>�"���u~s�e� �JÜB� �[�_��/�&-�m�M=���P��4vL���2�+ķ��&7&
�@�e%:�XQ�����p�hD ٲH�����USȮAJR���q�84�S]}�AO�p+vQ�v3T�?�"�b�X�߫� eS��h1����������.G_˛�����uj�8�%h@5j�����(cu�K
��8a��`R+����I�<��D/Z��Q5�V�fC�k��鑏���X�{^���LO�ʁ6��o'f^5&W��;�X��IS�eIg�B&2l�̅�W�۔4��PP�l�u���i36;_cc���	�P���X��IK��F�ݺ4��5l��w%އ�o�tk�eM
$Cp�TC2�r��i�  K~�4���������iP�t{UP`�i��ٮ;�$a�J~�p�>[�(�D�[�i��~��n�j�Q�d��#�4̈́.$bWoo��>����� ���l�+��/�GُV���<a���.3�����s%�i!x�&Ey���]�;��Hy6�����We� �1��5u������ԃ� �p��U4�?(6�H��%]tV������Ϥ��9<���s��T�N�k>8C/A����Q�nl���2�O�10�-*A�	aH#�X�rHgΗj$�q���+�􋎤���K4Xx�f����{��O!�0:6&�w�)���� ��ry���h\*8@_4����o�����;���԰�����xJ�?����}�n+�𡂨x:i�>mP���Xp<-��/���[��"��,��!x]�>����?��pr��MI�d�t?|C�6T��;����s���1�h���D��q�]��	����"�mʉ��W\�3���@B�u�Au��Gme�k���.V��=��Hwj���7֖�!�U�\ͼG�TBrZj��})��p}h�jN���-����s��W!ݸ�$l��Fp����;�~r��A�l樄2j�O]��M��;��'�t�~����΁� -&�3a�.�x�[Z��(�*u��Pj��������-���o�WJ���fޘS˲��9AK[�u�6#��=�긇}1n0g���V!De:2�y�6ǂm=,b�*�d]�bJ�e�M��1�p�����/g@�(�X�<����'�Ϸ>�|_id�x��H,Q�O�! �:G*6'���xB�u=����_�k��,�f&Qw�B�u&-�F������b4�pI@?�����e�����f�YbGk�-�+�OG �O�����YO;~OJt�� ���C,��f�@0���Y<̤܇��;_4�@F��m�̒]{�#�����&F�x��>�;M���[�Q���o�ټ�~Pw��@,/>(���Ԏ$��o��Y(!�<4�l�vj(d���n\�zm���$2d+~��%"_#(��< Y�σ����J" �o�7����Ǣ~SL��Cd<�� ɱᶵ��t������՛U =>�|R�_8�ֻ�qv���K�%���� }W�n��v��0����e�b��eK0a��"rW�UkCQ��]���$D�W?�Ə��=���[�4do�3�G2.? ��G�9�ٓH�������v��7��O��^]�!�DG�K�9\���I��E���vuk�,�q�Q��D�
��޳��w�C�N�~��Ѫu���$E}S��������$(us1'o|��֯��=�����$">$u���.#W#�W��ާ�!W+���E�m��H������$��!l���#�f�#�6�t�MU����Nm@e��>]�1���H��͞.n�a��hX�$v,���[� vl�:�-�aY�H�������t��]QFR��*j!N-5��)�)�O�[Bm�Sŀ�c��l�%{�R_�<w�e^�B�<dٍ� �}#���It\�Ӏ�Se�?�a�,�U���R�m�����d��3�U��p�Ͱ�!E�밀�^���#ml\���'��IlX`���_R�`�6���E>9.nz3E|��K�z�\��+��V</�0�(9ik���z����b�f���l�lb��GP����lexQe��w����1���u�ba�]D�ny�M/U�WH4x˷'p�����OgG��ڕ���귃D��_7�Aϛ.�eu�]z��'sf��Uj:���T
�����g����R��Æ����E��^��t�<H��:����;�#W6#��nՓ���T����v~D&J���%A�2�J�R��B�߷��;�!_í�=/0�꣜�1��iP�z{��wշ\��\�>���պ&��!ƙB����}�焋�ӕZp+�rM2W�%���;�o�����>Ԕ����!�����<9��K���`��b�-��?R�-��Ӿ����aK����-/1`�t�u��b�ҙ�)���~�cq���e�}T�y��)�P��N�}�ĉ@Ղ�]Y���~��&�iw�O��r}g���ϘLX����"�K�6���vP�JT�N��C�uw)����x�f�5�!��d�����(�p񦒾p�-|�4�`n�Բ�mq�=�Rpc�ˎs�[�I���3Z�#�w �����5��/a���J����-�HM,7v��@�hߝ8�q8��nm�+<55'O�<��OgSG|!��\��e�~��پ�#������-T��EQ�_�3�p�q�����Z10.u�E�jKz�`��c?~�J!���gm��Mz��Z���V��"Jy��]|�}��e��8,_��3]ru8C�h�Ѻ���6w�P���#� Y���1q^��]�϶m�n�9�]�ɶ�ʶ�lۜj�亲k�w?Ͻ��|��^{�c�\���Q����>�Ǐ�[��SS,21��"�e.쒓����.��"�\�W
���a���J�>��������摘H�3x��zW�r�+���S��AS����^C5�2)6ג�U�#�O8�o��^m{��`L?�o�!�"�Yx^��=oG~��71��ح�6Y�;Z�p���>
}:�j8-�:��뫌��~��n=�F�4Ɵ.�]z��iBY>�W�w-x���P�p��O�.�K����^���!�Խ�Pӕ��P�M2���
���D
���7�"�Ps�3����≧�y���� �=0k�}��3!�ϖ%?��|�l��-����y}�A���g�)�y�M��n�>�I�t6��ly=y]����� ���:��^}~>7t����Wn��ӛ)�b!���^�]�ђb�E���D�5x��Ǚ�E#Y.����~Hm!���VTR6R�_����v7ҰE�o�&;�Ҳ��5�����胃ݽ�����f!^�H5�(�ư�a�E�L�t����Ѽ���=�w�#�p��Qy��]̷�hF#�vX��wڷu	ⵓ$���q�`��*0O%ۑ]V~)�uN'8���G����*I�~>'
���D�6���*a�o[<���]2����x�ҁ�	�ib����O���5M��|`|��p0�t���ܮE�� �L��s�����in��=��x�s` ~���(5�kH�uȖ��>E����i�e��k;ˬ�Ί��~�t����i-�� 5�g�����I)rZE3�"R���BU��\o�rIkK������0�Æ�D��;T�}��@)œ3��滏���Հ�3"���6o�T	�65�7D�mѕ�1N^�����r��7���	�6\�\i���<,'c.l��}zW�3�M ��|��Um%�B�T'hh	*|ǜ@���e���t���;�H�m�O��j���[=�b/���i5x����d�o�C���?0�p��c^>�Te�qگ��z߃-���绷x�5u*��`�S/WO��
�(��=e��T'Ių~�r��k	�?|�]I��`�T��t#�i��C�Hҿ�.���|�P��r�p[�i���\���I��X|c��<���*�%~T�/6o�hg�o��7j�6�:4��V�t��xTNQe��91l���no�!�DE���y���ž���"`G_Դ\�H~!`�º\�le��8��(���M��bu�����X��Z��m�׫����*��b)N��i o�ט8�;}�Z��Ta�ȅܑ�M�˚=^���k
o���&�jt~@F.60���psp���Z��)L�r�J*��QB��s��Uy��x���84��;#[�0���v[-��"�3��!r]��0�6p����.G����6�\��C5a�Jz��� ��_�]�u�Ϙ`�Bu3b�c���6|���������уj r�������U��0ȏ{Ͽb�OqYWC�R�aTW���Q�r��Eh�0UaI|'��I�kb^���,r�c�Ш�>��ؼ���l�(�cK��ăᅀV�b�^;�\�E@ȎV�d �:��OMr_�<#���^h�� ��F{/� �:��v�	���A�qõL�>b�3�@D�-���n09���:�n�)NS�ˀc"������ p�W}j"�5e3с (�Z�E	(�f���f?t/��˕B�FrM�'�@=�-��j	���ibVFSs��<��jy\�d����_�͓6b����,5	-JUo��i�@#^�x�D3t�ɮ��`����}4���V�AnV\K���3aM����O� /IŃQ5�9EF͢�9U8� ��`n]����� � $7-��U�A�K-;��F��ș��vF��e��g��tE��i+�͵��I�4�L��{�[g[�UU,5p3@vv$��Z��dR�� �"]"�y��71��^�U1��N�´/_aU� �(���xT�z�-6�Eh�G�"��䌉E~n�F�����nr�>,
�9e���#rT�؇�R CM��p�Q,z�8K6O�yn���މ����p�{$��v�=��[^��t��p�Im����J�,������̋�^E���.6v�3��-<Je��v�̋� �5�_�C���^�y<�hn�p��4�5 �_k^��h�/�	C��*�Y�Ԛ�u�����	����09c�2Gr�U���0�l�ւ0��<�L�E��fN ����W��19Q�X��3w&L6l���C
��̼K���lO��qFF�)OJ8�W%ov%Z3ݣ��0��	''�Y�@�wH���O��Pz,�힯�O�Z��/}<}O)S�H4%9ʎ>!*
���/��%�)�^N:D��&���n�+�?,�a�H�tEI�Hg8[�E�.Y	�I���S�}@>�e�����^l>��1��v�4�!���?�,�D��1�o֎:Iu�ª5��X��d�dZ��mt�.E���q�|�b��ҡIu��4�PV%[�FL%��~�B��dŰm3�g$Ӂ}n"w/=������]6�ف�w��}&�v66�ߎ�Qe(���9���GM:�s�G�W�BP��1��_�>�ZY����i�^)��zO/'0�J*�<��q/�<�U��z8����N&�7^���}��*�Ϧ�r�B�רR��M#����d5\j6�!/���?����"�)�c��F�@�7)�i�^�?8�ߛLdRV$�1��g�S�0�S��S�f�q�2�o@SxpLז}pLi�<4 �1��h����a��"�η�\�x;�v>qDU���/�\��8g�ζq/Hr �HaW�"��Q� ���,��t�Aǽ�F��?����˾��W�=5�QK���>2 b����G���J#�>�y�ZE�=���q� a+�/O�$]�ᐍ�#�шD8�XO�.��wzsJ-��X��h�R1m:�G�ުU3fO��À6v)<��v��P��Ϻ�Ԭ��)���̺��F����jN^(���]w�3������.��a��TX5���Ȗ{:v�A�V:D�,�_K�9�/͖K�w����kRY��E�lğ�iq�=�!2���jh�&�\�u�&�ˡTemt,k�H���^��A:��h}�<��f�I�Hx�T86�H9022h5y�:X���Q@S��B�<�$�V�1����H��6�V�K��"���}ME���'w�Icl�����u�Co���c}�հ;u}4U��9�	�KB1���#X�A���������yJ-۽�m_6�ת��@I� :�༤��u����s2���?����H�pHf����Eg_�L��-S)]|��&L�jFziІi@���H������]:�t2�_���C���U���������jJ�	�D���.��o���et7����QP�]�O������k{��Pc+]MP����7�%��^�2X�ga�t��52��hn�#&��#�O�uJhI�ɘ��0荚{��-<|S�͗��t4f��҉aѶ�|||ȺuY�o��Te����GC�,�k�t���G�0��ƈ[9��9�i���\�/j5m��`�k+�RA&���I������g��svg?D�~��U�圧���e7��/��KZ=�n�9�b����g��_v~�Hr�[��<�.}�4�oh�q��a#���/�f����D�=ԨŤ�%Zz���q�� �x��D��RR��H2��0u�=[�G��}�>�X|�V��n�o�x��q.�QQNI������(6=fw_��<g�B,~�~n����r���X�?y�p�Q��OW�׌��vZSnA��Oظ�E0˂�<W�H<N|BQ�'E���2����Ip����E/�n@���)N�����mϲ�|E�O���V �<��l+h�,�A��v6�.�3�������^�{^��e��r�������r�ъ���)���{�"�.T:�d������:^u>/�;��������!���@ȃ`I�.�M��̯!�`�3̜�D��~�X�����z[,
%#Y���@K+��M���*����Ȗ�ߍ��!��|������E�S�Ik�**�.6���'.�Iw����H����ߎVv��f>�����	��7#⇙8�6����e�4v��MV(Sڹ������1�rM����Ch�	���f� ��u?T���љ��q��P퀿�dn��:�+`<q��y���^��%�D'Js~�[�����C<|RL&��Y��g��#�i��	lS��QѮ�8�2�R��W՚�QRK�I
t.�$/��_�kD��2���������Gz�w"h,�Yd��Ml{�~�m������㻓&��a1&�2:]��Kg��\����|zx�B��=/����E�&`����L[4I7o�o"���Β��ӆd�z�TŮ�P`�����o�:?�x��\���� ���F�â�i��VSd#(���4���`(�Ĳ�n����E�H�_��d��h�}�s��V�=�	Mr�������Wc���>Z��Q��܊=���;�l<}`�8ͻy*_�ߝ�@m� fw��T�â4��Ua"��DS�ŘI?1н���^��1ư�K���H<B,�5�BˠB*W���ԉc��"��b�疌Ge֠�,��87�׫��O��2�u!�#x�@-v�E3�������PL�|�%6���!����Lu���u�����OC#$97�>`����n\�{������#y����F=P����/���fq�%&ʖ�7�*�i����	�`�mΡO��7)�`����ƚZ�A�(�K2ݥ��W[ㅅ �BNT�m$&7*��T�+���2tZ�|I!B�սƥNL7����I�t*U�Z)��3�F���*%���I*#�g"~�<�U�L�Li��B���e/������RgK�ݾ3kC�)x߶�#O��1�v�4M��C\�c��I�?�R�/�"BX'�X�fg(3_��a>'�d���X� �6�r	�D\w"��e�����\��dp�U�zȰ[�NM��C)*V/m�\LT�Q���ah[VF�������v/�F�{���Ys�X#xX���O��Į�|7>���~��������<�\��}� #(
E�C�#�یB�2�|�3اM0��[��4H`K)b�i���h�~����{1�|�l���]���t�:��/�~ΝO�n^��r�R`���n��HWVq����D��%����~OX���!"��5���,�v�]��#&��8aģ�>��J�c�dV��{��������E�C �;CWk��y�$�} ���q�� C�����	�@`5�ul-Ev�r����^�~~�0�E��:���X�|}F�2PM���T����Z��`yr,]�@p���Ⱦ@���E��z$-&�M���`��b�QZ'fc�Z��Oֺ��}����dI����CzRc{��=�"#k�'�y�C
�O�"as�*��;o$���ҹuq����E��YQ%F٣#�WCHU^e�c:}���k��Q�1,�v��1�$����F���'Ȟ�Y�uLуy�-�٧��[�G'Nk6A�^%��S����J���s��Q�[oD�U'j� N�^(�8��ls�Ǎ[�>Qy,��$O�$����c��:�s���a�@7�z�}Q�����7��`��$?(�X��l�jd�yzT�D<X��#vJ(�缄�m�mP����4����ДO�nጮ'@�^���<#�Qӛ��+���wA4���V���Q�8�V}� tu���[2�Lp�>�Db�bm�*i�m�x��'TW�6��w5GৌO�Y|��߼�$�U�Ej���W��T/-E��90�E��3I�$��/ZȼQ��߿��z@=�cʊJ��P�r@Tݐ)Fں���<c��|ɢLeZbI�Q����L5lH�h�@�b�W��Q���h���SH�$�V�ߵA�P�i{���xV&�@P�n0���:9���E�*�q9܂��o�&npS���٨��A�D]e�`n�\N �����jӊ�ػ������܊ޯގ����e#ȷ�W�'�nH\�oЁI	p~ ��.�82�\>c�蜜�{VBO.���k��C��9���v�|�y8QCI*E�%zS-B�s'V;�9�t c<J������i��Fz�?�w(�#���,u�@�L����?ZF��ғ@�fZ���m9���6���w֌�A	cx�B�)�6i��TcE���)��a)��M��1�w��
G�i,%D������f܆K�H?��,���� ����vf�<�<�l���M��XZt�R=9w�}5�hc������tF,��c��iVrrX��X,�Jt������	�12~�C��������O�����W�Zs$�5��)d����3��4�T�:�y!��CT��y�Ŭ10Ğ&��V���?�U[�4MEL���z���ԅ��Kpo:�"�%A�7{L�E'
{q_d�JE�40;u ������N�yˆ���'|JOe��-��,�)�j�./,{~�#�2��{����hp��~�&K{`z�k��"�#&▗/U
dD�e����"֖RG�FIA��K��
�5��Sf��Qg��k�����Q�*V�KfR��3�!h�H�h��;�Ue�|Ȥ.5�$+����z�שb�2S;/6ȑ����V�΢�V�Q C������Q"�,��v�l�K�z�jSZ�}�',�4��w��̤��s�Z~h��`�x��xUl@�1�Z�o���1	�+=���D�a&��G����9u�i�lS"�.\G��A���;O�q�\s�� �hSYk�&\F��x�\�ۅKU��Ͳ�0J�p6we�b�[��������@�q�(d6���+JWX4�������"�j��oT����%�1P[G���ٵX�~o��i��N��t��]����(&Cs/$�9�� �`�2H��k$^������[~�	Z7kR=_S���A�اD�&���U��/��Hq�R��6��\uD�N���K��� ��G��(r-�K !u��^Jp�S���8�^(9)b��9��g���V�Db�*�hvaڴ{
�@���?�4�!�#�cC��6�e���i3�!^�l?HL^��N���b�����������aQ�[�y�x�a�pָ�qM��-��VU�#4��a����TF�#������dԲGV�
��8�45Gն��ёΗ�\*�w]���?�S���EB�8��{�HSTz�Ďx���V'���f=.c�.zx�h���{��0�f�3��dYL-!��в��q���5xz�abeB�Q�/��ot�c�lJ]��K R;�`��l�"Q��Q�iR��^�F��ox��!���\��îh�*3Β�������N��;��w����=c��$��XKӱ&s�O}�rR�ij��I��*������;��:��(a|FᤥaمCռ�ϥ��%����C��!<Y�"��W 9�*�������6�j����e=��W	!s-�b��aӁ�3n/ݠ�?1spMs?+��iy;ᆭ�x���ѽJt���d�D��St7��"g(��u�P���u�D�3/
�װ;�9�Nl�S�V ���&$��Ju3F�٤�Hı:^,�/�!"�]ec���QN`7�6dSA�Xzkҥ���T_�l��+ZX⸺Ei�z4�tҼ��,b&��3��%M��Cr�j#�=o����Xk�� �X�O9ݓ44=Yqd��ܐy�f����!Sq![
��gt�~�H	�^sʋ�S2����%C�s�Xfz�	opq�+�e���9�|e�Hrͼz�SgJVK�MNSenk	�: ����p*I-s5��7�����T�,����ϰoG
�;SQ� �hS���}������m������.:��qo2�\�f��_r��p���hSE����%��M�8w�L��:L�l ̟q�玲`�3]b7G��葐��������gz��Jh�;g��	^Ű��hJsv�yx�l1��(y�@*� �^ [�g$����f<K�����0X	W�l��f��&.C��O��������U�p)G}\M;Xnu/}�z�KV�v��n�����X�ۃ$`;,����F �I�d�f�u���eN������t��4F�x�Tdtꊼ�a���E��y]p&J	�����Fӥ�I�ƙ���o���R-d�����d˲I?`�W��B"f�Z�UEuZJ��b`E�q`����Y�9�V0�f�8�:�e'K�;*�Ϡr�����;�2+Y�$�i���j;b[�6���-B����${m2�u W55��Ȓ31XSX�6�go�n|^A��mc�*M��1��u#B�!l���P)�P5{>&�jD��;�r�tOS����98�Q	�@(������K~�VV�>v^��Qv|���U����чj�1�c�����������@2�٪� �he�B�;*xU,oγ��8����.A9�<�5+�f|�n��x���3��Oo*w7!�?�T�o1�x26/�.a�Qe�"Xj�,�2����Ұ��7S����#1+U3�Q�
���������O���h0�Q�!��B*@"C+q��fH�\�ޠ�8"I��'����g7�2)s�܆���1$Z�*�р\�[�$��u$�m5����I��.�"7~��X[�n����82�N^�$d��n��� @��;����tǅ�5�{�2C�� c+��!����ϤV=w�v�^w�E]ש%�Oc�� �����8�O�����[��`�����/�|�t.�s�Y�$ld��o����Of��t�]���[��9#����h�(�&��ǯ��ID�q���ڞ������$ն�bP>�
N�M:��nJ�b�5�g-{�Ki��Ќ�Y`�K�$}����^oo�u���m`o({'���6�#�t_EfC>���^ˈ;�);�o�G�Jd�WF3f�DS�\ᨘ�b��݈�ϡ�w>��Gh�}�L�5����l~} �������S�4�[<N�V��b6���fY�J�o��h������`�oz����ܺ:ɕ)/��}Ƴf'�>��C<\�mkrF�_?y?��#P�\�Vm�@	l~��B1��C�������{3���#�Ă�����F�+&����K%��
1��ծ����a�]�'M/�4�F�Ū�{U�r��@[�W�#o��1�X]<y��״hRX
t�2�޷��P[�a������a+~.4�ٴN������b7i�d���4(A�Jpb��ɦ�GXm��c�u���Z�Tb�P�v���P���bV�e������w���pT��˖1X+(M�OPD` �X]7:�.����In���ם�q���n��޾g?�Z���YFG��o�z��]y��&��)jA5Ԯ\n�D�T9�{��gvJ�Uf�d��9pyx�p�۶�Y�i�oBY��_�lL|���!]��~zO��*�<C�>��M%3�_��A��=6��\�X���$ּ����E��̕?��w�,{^����4ojo��$�tu��}숌B��GQC	x^�C�~Ba�`^������ݾ:�Cm�z�j&�B��|��wF���u(����_�CT�7s���N�q��	���:L�*�|���+g(����n��.v�k���f��E�6_�ʄ�-�4���W������BQ}E&~��#1-R�W��0�����K^D�}yk�XUͲ�㘙n�H�g�ICo�B��^�q�}���Nڂ���~��Q����ɧA}�R�O��饩x[L���h��:��7v2n�S4^�������q&Q��[������8Uv��Q*%� :����B�6+Ol7���6n�|����7��d�����uc͞�y��d�%��V��<7�@��K�G1xHa\��轅�Z�����VOT�o�N��ӣ����C�7�� Q���=�SEֺaaE����[ܖ���up,�hB�d�o�x����ȩ���F���S����b��9��[뽄����(�r���T`���މ�l�d�ݎ��v�2_�a|�]��ͬ����\�r;��D;vb�t�	_C��)�HBԓ�%8>�:�d�<ɋ���GX�'VK��5m��r�YG`�����GR�C	�]�D��������ż��ܔt�������zN.����?��N�oE��%���1Jvo�	~�f���CBگ�i��j8�V��F���\����:h�r%{����D�,�!ӗ�{$h��m�!t6�S\#�l��I+�"�8���ꆅ}�a(1i&�������b�.�T˨��6�|q�Q��'M��o6s#�~K�sH��<4�6 ��3�Zm��'�{h((*(�~�]S�[��`�S�t'�����Tr�7Q�m�/{
�Tƕ8���;\��d��� б/�|���8�\�3^��ωϐn��/y�������)�/ɔFιҝŞ&�y�G�:�[Hkb���Q�����*���#@�!
#�x�;:a�L�J����	�˽1�AS;S��a�{,)���p�P�8����E$��Կ�N�(~b���YL��}**��'���@y�9�����>b���W��{�T�O�a�/o�|�����U�~_�^���t��B�[����Y�_�PM�_�ⵦ�L���W�e�s��5�.;�tX���d5�����E�i��\�|�v���0���(6�j_��m
V�n*/^����T�{�W�ɑi7�ӓ�+,G~%��D��dEAN���YB�s�,�B(��;�R<M���=]��M��I˽t�Rג�a�	�I�������~�?��;8���R=�K8��;�*)��i(x��G���%��mWpG"�?;�ƭs��m�!�� ��y[�=c��j�qߓ� (�|Q�j�PSz-!��_V�{��l��L�p#�_	mb�	]��ܛ��y���U��z+j,r��ҫ���9�Xx�TC>#V$��4v�E;�Y�����jG�M�H�,f�2K!P.[H�O����`�^�.��v��u��a�K��۔BN�
%N�k��UQmt b�N�r�Y��	�Wt��O\�Y�����X)@.fA�{..��rcǋ��2�h��{>~�#V�ۗ� �XL�5�)Q�pK���'�������BN^ŊR��}��~B�Z���cE�9�BT�e����I�^k�@āO���	|�;��S�o�3�^���ȅ�p����*?��>hзgba1-L�Y@cHC���)�D��қ/3o�נ)o�\1,���ک(���Z�pB�?�1hln ��z����x ���]����Nʩl�@8���`�Ȇ�R��,	?uV������\M��0���涄��3?��#�!�~p-��]̔Ɋ3�d!� ����[�N'���W��j߽���˜���uU�'g�z��7����Y7���;�u!��|�mIh���KF�G�U��°�\t��?���)c�&7o���5V2�)�#(1XD����qO���ۑ&
�x����ۯ�f�d�kP�~+m��1Sp�0�Nf����Ȫ_��zF_ZQ[��{���XW�%O�Ws�7c�0!ճJ�z����-�N "-��K-����Gfn^�v�I��P��O(��n�~�j��z�R����7��H����YsT��M���W�bϩ)�aU��� o �/�X!��,��3���zh_���%+�b��)'�By0$o�nz����?�Ӳۻ�I�$(�4��״�F��c�;+H�KvK�����C8���r7!��/��� a�MGy���Kp[b�J�J1���w4tm�j�x�'�}{!��л�h������?���ʵ���{c��$oKNy����㕚jF�Z��������֤o�%Λ5����#�E�@���:C��/MN�a���(��i���)�_��L�~l��Fu�Fl���3��L��/z$�]tƻ`�f�no�_e���YZ���N�[�5G�0�G_��T����n+U/BH��*Z�}M����=-��P�B),	�γ�k[��,��R��@�-�K�m�9A��廫��g�)�"/�OM�)��]D�h/`D�3�K¡퓖I��-�¤��Zr_,�7�\�^����FL�����]`Rݶ�"�0�����������#�������gQ�~����Z�����-իN��>�'���ş��4�?�Z�8CK�qh��8���2�������	VFfd��^��#(د���n�S[�֠<�)��%��ʯ ��7k.��n�uV�*D�f�4���t���`ٕ�P�*�8�',��Y>��%�i�5��i0l���.����)i8+i,��%~�+^����+b�3�E.����&϶��!�@<�>oC���0sjQ�W�_���#4�NgqP7<R���2�X�(.+Ã ��Q�]w��{�=.F�f�9�0O�d�)���V��VP��y^�*����;D����b�&�U�˥RC���{���L�v}�#�؉�#������>��5�(!ձ�h|kBZ+�B���Ò��6�-�/�����KU2�Fa� �ʲ��JH�r���j`4��U8a:ucm�|�Q�V�U�;~a��<X��d�z�ǊI�S����v�����$�6,0�g�^IF���U�m�Vcd�/s%?�!��ǣK��3�H�hj��&�������^�K�n��P��#��c=O��_�L?=�yY!�5�\R�߳K�:��3H^�/0e�������������)e��+��&��F��Kh5�k����5���9���*n�^�r3��J��"�݌�����2�h����c��j@4�Id�ʶ��ݘ_g�� ��L]��)	�E7�L�r�xb6rX:��YΑ���}�Z	y,K��-Ag�^Ɛ��j%��4m��j�V�SSR@�p�/=��zʔ���cT�	}\a.h.N�����;�C����6HH9Ip�s����,Ӛ��ٙ`��P��J��8����}�o�����I�Jէ���a��Z$�ױ�W尪R�>J�*L@=��
;����z�6l�GO�o�j�d�F���mќTK�j2�Qa�����C���q8�j�QD�6���t�%m� �E������.s)A~a	�,��|;�Lu[�`_�Nt�-n����M�ߦ����>K@<*Jn�D����5�z��^��I���f�4VJ��A8.�(Z6��h�.m]���.��+%�2E�2[� ��+@&�M'KW���ת�v�[�|&%Pp�Qꭟ Y���#U��'�m�,'�K�9�"s�h�ι��mB��2�.��9�����V���u��:�F�{�#��O1�B�����}��&��<�j0��QB��i�2|�D��RV�9 !}U�A$[�&#�MN<���-�\�bS��E����Xʊn�w�Ag��C�|ki�zD�2\���9|K��D��T�h&!���D�:�-���Ss�IC�����eE�{i���Xg��,!�ա��Mlԥ|劬!O��>�\�}�|�e��e�\��Y6W.�B��-�͛��a�i���u�����M��m�P+�{�nSCm7�|q����g�6���H��n�Ek����K�Pj��:�Jܜ^�J9��d3��\WQ���1���ӆ�GGq�Y�gPU���R���p�J}���t�o1���"�Ϡ��GS��(l+��+���7�ZD��J�Ax�s.&�'=n��W�]�=��Jxa,�I�]-	.��!H���T�E �8�8tMl�������FZP��%�OI-�Ѿ��6��<���6�����ߙ�M�cz��1�wn(
Y���ԟ?kQ�2d=�m|�"^�zʪ��=~�%����!{�L�]n�a�U�ʥ��i����&�.�p�u�P��pH�\��(��I<5Ď�ns'���e��q���õPbP�T�n��fi����J4~����\���!�=��?�$욉��n2- �s�Yj ��`����0w�F�ֿ�&��dIO��ʆ*M2PTa�f�S`�K�;���&IB�ۅ�*�+��Wb��K��٫�`̔.�U,p��"԰s
�i�J:7���&�򘎛m���i���u検��6��2���o�;��*+��E�8SR�Ԧ-�Z��cųS�dG%�]��`�U���C�Dt���^�������>���$��~��|^��s�F�o=(۽����!�&�.*���"�R�h����;=�a����m�a(�@��q�TU؏=�z���F[o�&��o!�3��pl�Bt�����4��aywխкȔb��
�"�p��x�T ;ϙ����"�/&h�%O�Ϸ1'���<���<�A]�F�)��Kl� d"!.fZh]K��8vH��.�-og�n���UO[d��z��Q�Vq�֝�C*NUS��nRH�M��h�7� bu�,�E&W�^� o*���;�(��ZI]Pİ��|7|B�x���N��B�kVJ1o��G���b��wgT���wi���y��IW�B#v����5 Z�1F�Qͻ�;q� /I��#R�)҄j��ʗ�;�q�v_5�Ӿ	��8~�!P/������F��K�H�?uc�$��H��؟��5�m�F�Wܱ(��F�2�h&�H�{��Υ�jG�r '],���T?�e~bLe���YH��%����N�1o��mq�	����A+<�!.+r�a.:�ui�E
G,�������(����,O�S��P
�����<B�a���j*��O44s�n�pM8Կ&_
\��f�p%�2%����s^Q���:a4Z-�wLT�\�3������|_�Q�h�k��#K6F=�����u�|��{	��}Q�^z�G+
�8��a��m���VP�w(,dD����� �?�O2���5+��q	��∖��&�:�rRj�!�*��� B�O����|qd��Bp����SFt	Y��mgD>�H?�zޞTB�� 4#N�p�j�Փ���m��'wȷ�-����q�8�g��ׅ��^���<�0:0����G� �z�$>P�8��JS��o���^X��	0������w�> �U�j<Ɇ$�ݍEW�hj�����L5��Ǐ�bU�C�l�r�yο&#덢."0�����!jV�)m�.7��Y�B���[eu˩��!�
J�rX��w��������/8��(a����Aa��7�PG��	������pdr�G�'��6�5�����$a���1���$P�`�.gp?�Y̯?��,ĉI�(@���?6��)���=���^�H²�6*�VP�;��	?6���B$���n�w:Ntz������d���$�ip��]�ު���z��w�)��X�IA�m�0�ri-0�*�;���]��7��(��%)�0J��b1H��G2t��D�)x{7K��#}VQ�K���G���pL��MRii�I3�4��\]���N��v�я�A#��%����ƿ�u����߿+�'�հ%�&|�)�
%�bV�C�t1:�(m�ϟ�Yێ�;�ZU��D�v��5�ۅ�؈�"7tc�:';�r}oW2�
$:��	�,	L�E>3Ǖڷ^����\��O�C{�O�`�q<0�2�9�&^`J�仲t�(� ��:��oH[DH>�m��^�����jd�����z�˴H3|�vMɊu$���V��
Cm��AA�r�@_�'t�<�vv�"� �N]F~����GNP�����ˋ
 ����H��{�U���)��U'!o�O�����a�|�_@z�U~�R?%�Z>�xn�缉:�*���j��p��>�:�= ��Hw�$2�k�@�U��hQS`3��?x��ڿ�N�������p�Ǩr��f�������mߛ�|a�˅0��{$�\�@�_����wU�`�Z�rw���e�o/�	#�m�����3G���wޯ%����\�������TD�?��o���Y:�>���[W<��Ewfu����B�~�<���Q�:3�	�؍���<�sz�z�nX�0E�{	����(��l'b�pxu&���)epw����Sϕ@ޣ���yn�les��Az���*�V�*�No�wh�(��f��N�2����k�N�˷G�������e@����6�:��k7Ɋm۶mkŶm'+�m4l�4���h�h�6~���]���z��Ϝ$�ȁ퓎)4�EX�Θya�rc� �4�>�d���be
�_޻+)�'��q8���Pӗ-�Q��D���ŧkn%1Ӭ�0�_���8�֎]!^�#�ވ�-���YG*���l�3��o�X��Xh���Le�]�;��pN4G�M��-ۈ���+G8
��&%�	�j�W��l�C�_N�`���$�bn�3H����>��l:���o��b��"����,}X�aXԡ��(��"��2�6VeS2{g�-�+D�Ȫ��|�n�/%+ϫ܂Ą��B!�dq���b��Q�������_��(�%�胥�;}���H%e���
LR�Εp?������uK;�z��A��y
h��:N|�s�B�y�� �=s��~\���~� ��90v�6�:Sʊ�СR`�������W�V�n3Lc*�.�K�_m�Iv�������Q{�]�E\�ڌ���y�I������QE	���JU(=L�Ke=���g�{�G�{�7��d��� �0���yB͉0�/�dJ�+k�C���;����J�����7+�`3ZzW���J��k�Q%�h�t�;.��VT΀'�1��W��p��@�����s|~�|�?=��]�ӌ����4�;����"a�4�)7�ǅs��N���������ݕeDç\�,�^gJj`A{|��(�>���w�ǩ��"*�pF;�l�Y����n6�!χ��R�/2�� �p,�X��_�����]C(Ҿ�V��#��dW��__9�ɒ-I�ţ��q�K.�v'�E 2ڎ���u�@�T~%��5N�����k�dy�m}t������nH{�G���Ƕ�Mn����A>��	u�~��%����f�gK���
F����r���gՙ�f�}ø�,U�$����p(��#V�	�)#�9�ФNKW���GlZPu���qv�ו�^'��nPO5E�ۜ��u6�T�F�R�:�� ��(��qB��f�Q+�Z�j�;���{&Q�}�hQ�A^Z'�jk4 ,�1|���*�c� �1s
�dR�_�rv�������4��$�n���ir�!�=.�a��$A˓$A��<���w�w��=3	(��C�^�Hf�J�E�k�����L�,�4�Q��f^���Z�%PTs\fe����D���x�'�����o��<|�����v�wЉrsC�?a����ώ�4��⪼GP"����43���a��)Tb8%I�/m�,�M.�ܖ�rdt�܂��a�5�OZcN(��~�k���n�Z��A�e��e�̭��^0ci�c���u���H&@��9�m�:��Bq���ߘ"�2��K��	����ϑ!�@oUF�Na��̕2�����*#��ˢ#�6[O�` 3t�w��������$xV�� ��%�RE�{��$���)Z� q��M%�����d��/�{����c�>��Ha)*��o����|ʞG;B�Q���βtB�sH�%N�v� ��:����h����Rip�ө�m�H���,Uf�3 ;	Կٶ�R��A�W%�*�$[!Va��.�>���γ��B�@�	j��*L$e�jc~2WA#�R����H� ��z�(�����d�Us���o�g%b�E33i��,&]B�\������Ԫ��h�gr4�e��#�aưT��	�ҳ�;�m�Cg.d��ر����S�~���O�_�{8+�LvƌK�sz��¸8�+^�u���ӭ�'t�hC=��(�X���{u/w@��kf�ʄ=m��IF��y�x���Q���&D�
gP�C�4;h�*���^$�Y���/�1{K#�\*:��c)5�u%�IU{�_X�N<_{r�����1r#��������uƛbc��0Y�x��\��9��"7|�g��:ʨ2M7��Z˘M~�v5\$B�M�y��5��3;��s�(wێf�Q�Ԋց����e>c�|\���jR��.5�`�C䳒aC���'�'�{c��O�w5�.��B2l
�F,f%����wy�=[b�jX�͝B�g�ܘ"٣s�2Ft�[O�A*_�O1�U�i��Hp�a�'�&�ѧ��*��o�ۅهoMP��l�l3��`����7$.h��Q*^�;�i*���_w,���d
}4Hy�9c��db�&efB��Ӵx��z�5� ^ڶ.�� �D~�_*1���/�%Ƕh)A�^l�����̢T�O�}�+��O5�}�t򔻀-E�p��O���_�3�9�
*$t���eXB��S��S#p���tF1@�Pytʆ�:t5�=/J���sٱ�[G3�f[e���������J��2�@���H�b��/�W���F)w͇)���/5�6�s��'_в�'��~S��㊵��8J�#�ژ��98Dl���F��sZ�ۣ �V�ŀ]�������:jh<��K�D�ʺ� �EA���Β[넚�9h���
� 8Zg=6�?h��C~;���f5����3K^����!�+�c=�9rxN-ޠz��x)Er��~�+t(o�:�E%�oE���@&5^�!��������������/o�4�_��k����� ^dG"��Tb՚SP,�q@.��f�2|v"�n�À�C�v��R��̀M�-�l��󲄱�hݼ��	l5ٟa��`����g�S�3�
#?�9����@��8�G�&�mѥ��,͌w�Rl�bl!��!Uj�(��t��G�G�'�d��ĝ� γYH8M��N�%)����]�b�ᵈ�Ϙ��qwI�(J�@Z�^�����|w�����m$���t~?��E�R���8��;����úM��n\å��7`jX�eO8C��� ~;;R|6	�,~����Ǡ+P@|��xM`}�X_M���9<�[�c������Sd����M �ݠy��^>)Epa��y6�,��6�Np.�t�a�M�
�a�3���,Qz�RM��`gױD\m?��XS��Qn0}�g�J>?G0.S��h�<�L�9�`�D��	s���0ϣ.��E5��x櫶]��T3��/�	(2Z
�:I��x.�f�l_i�}�F���L�Q�����Z���|s�^��!�ߞ�8�L��SF'�����Ʒ�=��v�:�������n�&�x�:�(�P����������|AgV��a񶢸�E����|��|wi�����~mŁ�g�8M�ā�{!,bu:8j�	b�Z��scȹu����i��z4�e4&5O�_���D�	��]��̈Lˬ�����wL+���(!�ݰ��οj�c�[Z�鑌���T���W��7J��FWn��j��ov��R��Vؓ�Seh��>�W�۴��'	�ژ!���g����ЮP��ڛېO�*#�˗���1\���[�%H���ˋ�f��Ȭ��=�������E	�s4���%�\'�Ϩ}�Q.�=:� 
��\Ku*��r�$��M|-�����/Y��+���
���{��P���N����'΃�K�X,*G������E��ۨ��)��t����z��e�NB`�硎쫚,v�C뺊��M��XMH�m�L�pdh�N�Б���'G�ʅ *%�	�#�W믔��	�w��곫6�f�X�����k���%��f�m�*�r~E�sWV���s�1�H{����z����͘<���l���ŔׇjFu��i�fL�`�\"�˸���O�G"��Ɇ.��������R��U�� �������@�=�#�]��#�wG��1H���^�˧�G�����u�"O��$XU$dHc��Х�����I�-�N}���X=���Tqpwofvv��%6{�����I0��쐆`1�����t����^�W咍��Z0�~�[�e�`��8'>R���%K�!�׭o��R��}��зY��]�<}������*B�<]!�g�_I2�KU�K�gKwl���b�-�W:O������{����d��H��}���o�4+{��^��b������Ju����|�׾N�u�Q�3�5\?���,JA��b�%�!7R�	Rn�~JDc��}	����ia$��Ӳ�:����[ai�"Py��I��i���`Qʔ�e5c�@�n���w�Z�l�1�P��ch���;��= 3��T��:s�3���W���7�H�m͑(��Q��U�Hȶ�hQ����s}��x&�`�+g�W�8'���W���2p�Ce��� c�LQ��O~x��R��ےGޒ�5����ʭ�����H�8���]�0�_U������;ib�&�U�	�3N��'3p�]Y��4#��'�]�7X��-�^Z׿�/U8�.Kt��$y�������K]v2I�]R6Z���� ����C4z��o9���{�u4J��X/�v9ú�y��g @o�z��dA}�8M:�g�� qu  7��-d�J$HPۅ������(6�UXz�����}ރ�350J��Ν�#�5~�^��o(i��u�k��
��?5��Ώ�Ck�rک�y-xX�4	R9��	8�x�֙u���H��lZIRe�G��)�}1��W���v���Y����MΔ"?U�U������C �k�pY4��*)�9��6�'�Ͻ�8E~����ҿ��4T�Ӗ��zc�%4��!"~
6�;�h[�<!�u���0#��.�G��-�z&Y��r-��~���ܶ�Y=�����jp���I {h�fe��U��8_�s�X�a�}2�f�&~Uq�Q�zh���~�r�eA���/T3��P 2�m�G|]�ꍯh��Ɛ|>; ��6+�i�-�q��Ġ
�B��S"�}j���3<g�w����!�G�q&�D�Ue��dqh��32�l[�2��~��B�b� ౨fA�.��Ӧhȴ?�U4ҝ�$e�x���d�n0�6�Lk)��ˁs��/�kK6a���B���^W���w�R���Y��yq�}�WM�y:V2���ZF7`Au����^u��EgR�rQ.k���_���*�wV�["P�ҿ'�J��5�W�&��~�e�M�������O�v��B҈�vd�Y'��t�ո���!���@ԙ�'�����n��s��7�s>��'�����T
�B���Tx��dRqz��	oD�� ;o�Q�a5d^˱�d�Z(q��_󆻩��S�xH�
�y����Ņ�#,����U�Y���:�!�y��*���u�Ag�W�G�W��x��J��|\�W*�)�.Ϡ�� b�a��1�"���nw#����,��jìۄ}�r�(��Y�x�o���jm�<ŏi�l[�Oޞ}�o���N�W�V�4ƌE�SG-�l�v�����4�<)��>�@��h��[�����*�eX��*Xw�
f���!�W
Զ�ԙ+�^�>ܨ{��P��u"th�?��	;G���ic�i"Y86Q�@�kl��Vy�[���%q�
*xJ9�CN�n���'��+Ͳ皂b�wc�/�I�5���i�{�{�)���\�jc\MhEK��VT6w�mSF�c���I�G���U�1�c�vT�<�1`}-�rf�b�4��Zܖ���O�$,�lW���L6l`%B��� �.}�kA�c7ɜL׾*4j�X]�j��B_����x*�h���S]�����~$cQ0�� .�o���l�z8]�.�+P5�.IU���]��a5��&�2��ৼ%�q��-�0���̉��
zR��l,z��5U�e�RP6�˼~����5J�܅_"��=I/� �#�P��6Ϫ�K[�7��e�)P���2u' �X��_�G�f�I�aSعlh����!bm����LW�b�g͍p�ù�'��Q�kt��oF9+N�$�(�A�0���;qr�B�y[�Ԓ��.�Y'������Z�*<Js>d�y���d	��`[��'�P���(��wBM�>w��M��[�6<!9��V��ѕ���q0ɏ��'o�2���Z�l�U6��������j�*��P��q�͖��z3-pX|j�=�օ���;,������^�-��)�-&r U ji��$]�^�%$�Z�{���A0�~��Z�B>��\�/u��3���^��MQ��д�;ܘ?U�ȼ f�J�^
u��Rr�{�s&E:j�9�\�;���G�P�ui����X
�	3���8"�����+�|J��G	he�f�/��z,�UX@ �K@bڽ�`��,6�j!�>�mP�w��I�׼~���A��}�$�T�h���_��d%��S�a����� �Qϳ�]F[�/s}�)~Y�1��c���T#��Ā�P��*���h����,�J�z�غ�4�;p^D�<��ʾ�Ok���H��?(�[6lC�d	�y�$э���ѱ|�(�
ŦRs�y&�9���g)��m�*��l\L�]bο��H����]�V$����vt/���G�w� ��\��{�WY��O%���!��ɵ�sU�,Z��%gY�@�0�577�1 ���Xq
9���2O�-��m<4��� �4ŕ�����1֗�}D��P�G�ry�f;sZ-0��ƴ����ܗ�w�8�+%�.	`�Bw�˽fE�~�u����a[0J
}����ta}��m%�C�8� TG4����a�7�SD�(���$��e���eSc�r�VJ�7�Jo����ë� "B�"�'�"2���Ӳ�"�%∃�j��7���M�e4����e�7l��m��G�-5��ݰ���tk	��G�E�A;6V�yI�*}4������t�g��M�VOi�}���Bu�'Ն�q��'�]���H 7���Ӓ��hd��煝#g���y�T>{��&���e�ʁ�J1�{i̓�,v�b�6n>GO�����ⰱ_>����S��g��դ�Z;]ۉ�S#�}�~����O���G�˅	� �:�(LQ���+jU���>�-k3}׮%/�M7G��4��7�d���D�D�aת����(L�S���Hѻi���^X�҇�I$��]J�5J��f%�m�JO]�e�U�� �d���n�̱N�s��֝;R����M/�F�hP����L�i2�{���6_�S�Y1cP5�_��P�[�eZkTlxt��V"�_�:������1e14���IVO+��?��x�i���P�}��B���p+�{�璿i-$w�5~2�؇$���K
��:K��.E
���xdBt¸�K�)�ߺ#ޙ�ɚ�����e.�%��^�~���mǵ��G�m�S�آ���6���'��C�Z���	���e�EP��2,�x�}|ۊ�p�C��'�[鷐��K���K"�b~/���b=ʯRl421�P*L�*���	�u�ɫ���ޙ��L(D<S�m����ڑ�˾��n��S� ��ƀ�{��	�f��U��K�O�K_��X��(�2[\�v�]4��MN8���;�/������(iiϒ<iL�'$���MU:��J g.W����{5��7�}y�_f�˾]�Ӻ"&�>���r�O2��~%�jH¤���s���3Y�:����9!\4��7��S�{��)�f�]r���4c�s ØD��n�d��H%F���j�t
ذ���&�Qx=�*���~M�l�h�V�3~	�y�M�a�p26�i�虞D!l���O�8�᱔���0���]m��1�ER�BMy�����dǝen�$���N����86�¤�hؾ����2�8��|LA�h�C�%�M�3H�L%�m�6r��[��e�Pwӛ�Ӌ����Y]�o�K�hs�37�����M��)Ц�2)��슋�+�n���|�m�c�u��;���)@��"dbK�T|�~`��+<m�����,��A���j�Fk�{�(��z��U*�;�1��"u����H�}
1G��͠������͂We�����ڱ_�9;��@�dk��z��;��uak��Y��ŕ���:�f�|!g&��[@�M���S�S�~$6k�2��ƌ�����m�>�a#��TR�[�8j7�.`�RI�gAo��[��޸�����.,хqY�~��bΉ̛-A�e4U*��_���R,Y�9�+=Gs0����'�+"N���¨�~J��9�X�,Eyz�S(ڨ��zb)m��ʸ���]�ojf&.�9s����I�0P�d4��۰Ş�}�E��U�����7c�􊳿�_��6u ��حW��Ȋ$�*~~xSt�����g�NN*̗�7^��K;�;�9KY)F�"���#��X��*;A�����B,�+��z��[!�`A���kp6~:(�;��c��(Ǹ�iè�k�����k�l���V�Y$���{�<�|u����=E_�GI1e�kT�A+ͱ]A7�7�1����`�F�/�c�3�ryd��V?�P�˞��˴��l���������';t��7��5����9�p��6��hȲu8~����$3��2�#��t��w�6�1��.�y��oʤW���Α�0Z))���]B~�C����TL��M�*�lvv�6�ڏ��z!1&f%�Լr&�&��lGξ��^O����jA����0�VBx��آ-�rX��]�((wt�3L�H��I�Q��~Յ��^�w�x`�n\�{��W� �&Q��4�F��<�[�y���F���!��
�5�3�
��Kq���R�An�إ*���X�{�"�9*�<��eA��e\�i�l��룛c�`��Q@�r؊��˵RG�sp�ø�&i0
�)��y��^�I"b�3��h:��4�\z�V�����!v&�j�Q��ԑ)A��+�t؇������|����\�R}�`�񟶤}�g���a���F�k��$�9	�,�Cv��C�t��V���L�nN�̘S����M�%� ���yxS��D���_F��}�퉴�哾�c�c����-�j@����f4RX��H��9�)wl9�=$"�E���}^`��MW��[,�R�_��"H�PV��@��JR��^�!��4�k�g����a��F�q�i'��78Ǣ��c���ስ�|�eZ���#^��8�^ 5�((J�!ٓ%ޓG�^q�SP̐r̸y��A�=�r�7����{`���D�K��3[�����T�W0�K)��p��y����'����	h����΋�#�3P��EL�K�R���8��6Q����@��Ӄ���ӫ�ߥS;5�K=n�r�G���9�5�P-}�zpk�V�S���O��yg0-�D�!x}�{����S,�ģ�������jx~:��>����q6��d�F��Ń�Q���]��x�h�U�~[�-��>�5��2؎
ݢ~�4�i�f�kx&x���s��\)}%4�>j��Af�W�zT�!�4��,O����!�q�a��e`�3aVh�	���HO���kbi'��K5�vX6%�4�Ă�bʗ��+g�]�8S��Y�v��$z�E�:�~��m��`?08�,*�x�]6[�ȩ��N�H�9O�J:�s�c�*ǌ�!�RːxRSy�G������'
�C�@�A��@��G�j�!
3=Wg�o��@{M���R�s��7�d+��6�&8A\��?4rѤ��$]�����$=�-5K�ɋ9s��xo`�w�}v4U���'������Vg_���*.�;�Px�ѭT�j��L��csU����X19}���C�$�ome��t�ǋ��j�N�������T没w��7Rߥ�a���w��3�i2�N�͙�N~�|Z���X!;��C���r���)J���Ym�Br��
�rOD���3 Y��!���5����L�����2�z�AP��FT���F��T8P�,��Z��w�M��:
D'�ڝk��h+�$Q�g:�+D��CK�ER-�0du)l�1:+���WEAZ{|~֐��ªO�)@�&�-������蓕�=,d�2%*�
j(��s3<$��������w��ʸ.}xѷt�0��f�h��hQ�jY��QL>_[R����3��w��b3Q�:�xzc,f�*�b���Oន#wo�ڀ[��4�t�Y[v$צ�6�� ���(r�2�����(��^I��[�چ^�[Y�_��ﲺQ� �H���r�]BH��%������bv�%إFd6xs�>ͳ����0ߦ��MxF�:,cQ�>�ے� �x��9q���So�;�=w���|j�%�����Z�7bA�d�W�H&bNl�&��S.�x�Lyا| �G�l�W�3c�����Q�eB�
ݚn�_�n����@A@y��h�ԗ,V�����_��|�@���8�s���h�^%����<���Y��U*���{9q����0+KCUQ�(��c�;��!�I����/B������t�z�8�u�$�ON�z�j)��4ѐ%����)%�zB�j;!b�ݖk�/�{^9z}s��%~x�t}�
{k&â�i!0D{��,UĕK!_0V�o��:��?�f;�o�.*�nY[`�ĩ����0	�W߲`{_�����}��/{!|�H�_\Ȥg���t���D����ɼ.ڙc4`��>�q�t�ܸ��w�Iƛ����>ȱ�Mj���K�?'츛��c��b��%s��N�`^^Jy��f�c-�:�$o�cg*`s"��zm���Z$��*���Y����j��wAǓ��W�=�L?�&q��.��D��Ȱ���a��]���1�x��k�J���FEɹ��-R�b����S)�Ck�5fvZ�c�Me���4���v�{��k����a!���,eU*��-�G"��r�TM��5X�~,w��p���@|eG��[X[��X��e�5��u+�|�i����ܗ��c��:�Pv����D���]�����Y*�[�Nve�C�q�[�c�h�"���9�m]�]�#bl�G�VL�����]��	�R1�66��8I�(����(6�-N��Ro���������r�`ށ	����Bl	�b�I�E_M�^^��ԏ��٠V�� +����#�5D��_U��D�G�����i.�i��S26�7Sg��nJ^���Ba*g6-5_�Dbz�
t�'	���h���D�L�����q�����0�/�}g{N�OZ����T0/na��K����;��㧷��M�)O�@�蕯�}o.�0��B�g��:J��&�+�FE6<��%0T?�6�DG�(��@\i�VY��/<��*of�S<I�=�.�<&�z�L�g.[���+d�'��>%���Q�>�&�'�����"�}Ǯ�y��h���9��*���1AB���.�!�[_r�y94��AWo�����������)_�Ϛ�6O��rB�p���i�o��d;��X	,,l�n�.P��i��1�5��j%L6H��uX�@MɈ
��@�W|l����E��cs�4��:5c�)pU��`n��x�p�G0�ZTۤL��ж*-�����9T�b,~� x���\������~���7�M�Ȧ���DP(g����
�bQ�~��,d��Q�Z�z���(1Ba�NM�v>��%"Cl�2,���iX&&��X��D&�v&�l��<q8-��v�+_����y�gB�J��D$ )��-�t8E!� �VA m�Vb�d:�D�O s5���A '��T$������\8FSX�%d?�H��F<�1��� \ܛ�vA�n"f���~)�Z�v������3��d��@���UÂY^�����Ґ�sT�
�\�ղ�*�(9��bk<�-hٮwkrk�^�{y�����lz�h
�'��U���W�&����?��/p�ʴnM��+7����oMpI�oU9����3CH5x�M�L�,�\�ј��K!�s��I��j��|���_	`�=I���HB�Lu�M�{\��UHc��fד������'`��(�y�F˨�g6�D�����Y��|�d_ϕmhD}��PPD�i�h�%`��FM7_�^����V	��t�;V8�aĴHFii �4IU()�����B:Ү�IoL��QK��<R����T�%2	�
�Whe~Ŀ���f `{6Cvf�RK:&XS�?��1�䕑{RR���mH�����rB���^4�����c�C�Ao>8,�;�0���I�GS����e�ԛ���X��"Kc`�ŠD�_X'��@�Tg߮�qg���`Ei�́��4�+^����s��A:bk�A�<C��4j8�[��K�N�3�����Q���?ym����<��f|9��C�����T=��⿙ jw�Չ��s4m�2�-�IF������خo�jz�]�G`�Q�Ą'`k��*(K��L�%��|ɆV���5!��u��KJ��e2@���P�Yנ�T{(����o1�r�B+����� ֊���Hڻ�2�K���*t�k��\��$ߗ���w�<DPK�<�4����#a4�i
�D���$�(��+�C)"� ǜ�K�\t*9F�=�Y�C>�B�G�[�`�7���7��{��!m� T.�</D�����=_�	>���@V��v"u'_�F�����-y���w�<���3�S���,6>6�Ўx��AQ<�Q����-JIN���3G}���8ѮD��@��u��XLC_9�W8�e!x�
@@o�l��4�C�T�*l�	��ST���W1X�|�ih���ѝ��qӹ��δ�P���	2��$"��[��T�3 ��:�JN�ȡ�ޑ��pD2���'@�YG��Z�L��4e�W='�sh6D'}�
qq6d�Qe���p�P@��3�U?��/"a�gM�d���O��3^��g���o��~���2��%)������$��
m�f�etFal�|J�!��YKU��ŝ�]\��L���-��8Ҁł�|6�8�z�D��(��!Y��Hk�nEL�,�h�L@=��\hr�5}{��*���_���8�|��q����9?JꊬVe��$�[Juǁ��W���r���Qq����_��|������³�ζ*��aU����A��-�l����:K4F�b��\M*srbR"+� C�"��s]���+���S�*�P���ׯဝ`��> rK.6�9�|��IAstT
!$�].��\�_��L*Mvz��9��.���Y�j_W%�V��z��ï������� �/�(�8b��p�Uc\��	_��ӦQ/�+�rYl���5�Z�㛁�9/�óe�4�lY����&����H�l�A~ڠ7�W�>��5C!�zh� KF<<�k���v�$��k��2�z�O����C!=�o8|�c�ͫd���zKa٬|[Te��W����Ju8����uF�Oh�B.���nbE?83p�M�H�����nF�lqf�ܼi$�:4�����?/}��&��
��"���9趘��q���G7��k��s��R7�p;�qO�Gc�^^� EɹiK�\s��@+�f���O/S��^f��M�Y�U�oM��V�>�� ��_H!�H�Ǳn!�b�f./�l��1��>]�b�HF=��oC���l�/���7C��~�VM,�K�>�:M��7`��	e�	��v[�� ؏��0��wa@5_�bN����\i����)�X�"�R�Q:^�{!�I��<V�FA���m�v�M� ��\�#�0��PJꒋ���B�C������M�c�h����^Pm�����q��`;i�����]ƴ��?�fj������{�=�{�����I䙶xb��S~�s֋2Q�d���)9���l�I�@%�DW��n�=`R�jl�F���?*RJ����3$�:[�CC,[�}M9��.��4��?�<�?]�_��7��i�#����b^�.ڗp?A�wD��}��m�Cd(_b�T�%^R-c��D zQ3�#�l�K�sB���}���F�|�	!���8������U�|x��!ߥK���d%!)�ũ���4��C�~�^��?E,9�.��F����z��u��?��g��Ȝ�� ��_�ڝfa?!���f�h�9��\5`n�B�q���)���Z����,$=��(�?��"V���F�e�,�݌�' �y��oR��nN��w7i��T��H[�ۥnqqqD��E�x��,6*�Qux���2\�u�k�RL$z��A-�Y2r�u�˷����M]
*F�ͧ�`�Yؓg=�'vd�r`��V������������e�{фTؗ��n[��W1��Ѵ�]�����r�匼�UD>�dN�T����`�&/�C��ˬ-s�ȼ��"G��-Ƣ���E�s�*f����O\�5H��K�OFn];રtA�֏
�W��$E���\�_�*6�+�9=����Ջ�A|_�<�}?{^�G�K�Am&����"����I�Eʳ֘f�=t)$�b�w��rt��k�����<�H����0�:[�����1��>Ԯ���^������O*dN)��y����՚R�߃���eU��V�c$�� գ�9H�U|G��褂��>ٝL_�R@��|e�L�~y�s_�6�}�--�_LZ�� l������ 'H�J'�N2E"��jY��m|��;h��.��Nޯ�-�0g��d�������S_�dM�xE��۱� �|\hg�[hlrs�)�x�:�|,���l�X_�T4���Jc :+���l��=6���[����3"Rڮv*i���'��1�p�)u��,K�B��bq��ݲ]����W;"�!~��ǃ�3Κ���R��H7���쾧�5�5�� X@�5`t�C?�k�􄅦�Z*&h6�L���꺩��Hm�|�q��qe~�L����M�U��@Iy&"+���p/NP���R4��G�Np����l<Z߉Wd���bO�[#�*���So��G�-@�_�j(vd:�h�]Ӑ8��~���|~���լ�4�#|=5Ov5<ݻ܋�_���"���3���5D~�nt��^R��ȼ�A=/P��/ה�!�.�z����a�r���eYM|J^o>��������G`�w�~�{JT�i��\�#��(�r?�ʢy�����P:g��?��h�Rx<!��b����s:3#'zK�S6ӺT�7~<���\��'���,��ٷ�[ĺ�t��@�1�`�5I�x�2~�3P��L�K��q��d�>���]y�Z���5��6�_.�`HS�������Cݗ�E7R�S%���^z���K�`�#����E��.�*G�Y7,�6f_eB(��������o�YQ����m^����k`aN*/�~�o�x��{�5���򋍡�
*4��[=��C��>�O!�.���A/]U�kl��h�����e�@_>w4ի�#_x���Y����PɔIjKXX���+�?�D�[Os���b�d����QF�-!��P"ɡY��Ҵ�.��.�Yp{�n4[ِv�l�^M�()�"ֳH��|Sy./����C}�R�^�H����{PI��ŵy��;I��rH,�͈��r=Q��_������=�U*��	����c�D�[
�ݴ3o�H+�w��$_�Q =U����j�A�G�֤�>?Yt��Rnj�	�-�q�SR2��Q�v  ���b.��n�ަR�^�#��s�+�_L��Y�xf�&G�#T0K���rX�L�-����J���MV��x���]�@�(��5��:�h�[轍u�y�+lD��憒����"�)~�a�s�ݞ�� e�CA�<�eW	#'_��܍����B��J<r���C�N�5+eE<�E�Ҵ�E����cS�`0ze�Tt�������@�6�/�zs�3�+�V���jY⼣�VdX�m�o�٢�0=��.���/�gɮP�t�羄��4�º0�<Q����^Ss�W�
K&w�:����k��IG��o��>�0���י�k�5zR�Q�G�#��[Q����]�0\���h�ڣ��e�MBa���N|=r;��E��d|��'G���;��Ɣ��_��n�5f�a�e�ɢ� �������Ɔd����fL:H*�M��p=c���:+Gˠ�K&j����� 7�	}��7�gs}͍tp�	ʒ�^}��%Н~�V���*Y6�0Q�M��bn��UF�A�X���8�����f�1��y��(U\��}/�b[�WŠ���^�A��D��[b۽��� �#�l���|�J<7;�:	�|+�o���<~�Ѩ�"O���E��?IN�Š���_��x��7�=1���ո�"?��Hj�� �n��W#r�&ux�\'r��|���DM�PL1��M�,��>�|S)SO�@�~� �~��>���k��b�V	����ge���	4� �Pw"RY,�^�l�x��Ǥ;�W��K�۶�tl۶mg�vǶ�ctl�c�۞ss_��Z���/;�%J �L'��_}0@_�L��լ��i��� ���I������VX��~�L�B%/��-m��m�V�蠻�A���>��3����'�T"L�0d.�;��	.��"��qH�hy��@nwM1A+�9�J�ǚ�ϲM�Ԙ�m�jRh�=�Dr#&(ʛǛfׁDz*�.�\�� ٞv��p>�nn�P���������m���G��"�j������7h�%����p]���)��'��|%���N���G%�6��r��e�(mgYt7���k%��Yt	�R�em��ĞYB��?Op�Ç�f��lN����m�1�#�'��ǷU�8�e,S� �A:��yG]$��m�Ir��a9�_�;ȗ��<T��ƕ�VVsٍ��d�Sd0L\#�>H%F#ċ��Wt��'�����W��Ǆ�6h4-���A|$c��b!�+�Mo���]X�,�u�z�꽺�� � �����N�xp�����	<P��k-,��y�� 6+O�Y+u�oV|*ښ6��I�%���'ЫwT���^R"5C^��󧊕��a��u:�5�to
�"of}�PZ7l�.���U�Z�*  �G���^&z�
�#ou}�2Y5	p�v=�1��З1]n1�ڐ�cz?�s�G�nw�>��1�/�Cmt�$�c��$J�*W�#��ê���3��Qq���#$���� {z N�� ^��'ր�K#L�ÛHs�2� |��7��]�E�0fz�Y�!e�~���������PpO� b�̙޿%���M�����M��6�Y��ﹿ�:�^<ij��TL��lQ)��X29�x���S]�2	�{I<��%���ٮ�C~*�]S���Z����C�m$!a}���R%8\�(�j�c �e�e�*,��� iX8���-�y�*��.��h�@�W��Q��L��gQ�(��NV���8Wvȫ�l*V<����2,z�g���B]ڤ^��$�-`�7��U��i�����֬v��5(
eM�,5��O C���Xo��/d�B�S�p��r��������5�عZoY�$p�/��?�3������l�$8țQ�mV����ؤ�*����Exp}-L������8�p�@h�a!9���y��{�Sr?In�`UA�ZLߔ�M����*e���,��D>�,�*'F�D��K��	΢�����o�q�Z��SC��|�f� ;�U[�JcN��S���Mឣ-���B��Yފh�*o�A��G�)�_��Q2U��Ɇ����G�<l C������8#Piv���!q)�ܑ���|
�����t�Q7~�>�>�!�aA7_6�@�:��2��8�5��S��������un��Cum)����A������M�U���!��WNIiM�/�OY̖��Щߎ8���h��q�c?<nUG��8'I5d�Xp��s���s����^�����>��8!朞���7Iv�M��8��V^�ʉ5�B>(#x�![�CQX8\�{����)�x�4@k�_>u�e�||B�����.p��'^n$��[�|4ۇ�*�pr�(W��G`�vu�?�	�������9�G]�[�D(�S!���9�x� �2���N-�
��w��:�&�Or�k�b��)֣�o�a+ r�mQ�t(B�a�k��,���6���0�0ht����@�c��K���ߩ�|��	������S,9�.#�Y74E$��ȴAUרMxU�����pˎ���V�g� sn?)���[�!;�I1"X�/ʑ!Ũ(w��əz[A9ѥ�T�A1�C�j����,u��yE�=Gl[�V]�t���j+N?�ht.���i[띢�"y�v�5e�t��������G��v�	��DDﮖ��fͺ0լ��&����z����1�y��q������w����1����3!p+m4�c���x/���X�f5�d] �=��I���<@Y�W�O�����ϧ��A���+��0�9����Z��zA��z�J� C,������k{t�m���V�bv��:���{h�:pe����'d��5����b����>2�2{@\�L=�],�6ԍt�]�T���2��u�*`R���ܱ���>��Px���?�y�f��f�Xe��g���郋��5�-���ҧsZ�H�E��N��AHw-9� K�Uh�H���&Em�d�q�y�c`��9MW ?{ gX� j<������4[7�Az���x�<U-�Y�5��]���u7J�]����s[bu���q���[L.��E��P0,�����𙰼1��0$�����
KW��, l�쎴�_=�F%��=K	��?n�_������,YdFD�N��^��6��
�>ZN���7k�NH�!��dVA��V��"q���7��m��F\.=�Yb�I�a���@[	�$f�@�����1���mߞ_�[fX8��ͻ���w7��~v� ��fMr\���U/Q8��q��d�c�) ��������iZ��}I+��9��D,ZP#[}��,���X+:�c#B>:[8�iC��ڦ����c(})�V�{�4�*���~�~YG�@��u�\����s�d6��� ���0x�	]��ڒ�ttuZz��=c�$ǴwJ��+�x��~��8ve��9�����D�|�1��5����Ž� ���LlU�0#h��Yuj�e��F���E�ȡ\��f��[�IX��w2̱ˠC�k?@�t�Ū��ڂvk�(�c�݉O�\�t�C�3y͔t��	�R!���F���ƭV#\�)ǆ�&�G0��������0M2�hkپ�>��݊2���`�TC���w��߶��R$������	�­
�f]��w0�9��JYuωo�͝��ͺ�� �w"!�Y��ĥc��{��f|�F��e�k���£Ða���ϐt���fީ?8� q��g��&OmI|���~�%�c��������a�����+�1Λǀ��[a���x?�X�?�B�J-S�i�#���"�.���#{�ѥ�n����o���u&�RdvZ�B���zY-���c_�7!��_����Q�81���p"v��(�aINU�l�7"�)u�mtY�B�����c������?��C��$3�M���g���I(��U��%��� o�����~���G���?�p�=S�|�A��ֈj�d��O���J⹧�)����u��Z�(���]a�*O"�]�/Z���梨@��ٻ<������T�-,^,�'Sw.���]��]�1������&��ݫmC-����{jW����n9���z�z���U�H���KsR�c�ߌ [����Z��+���p���;&+V���u���o�]7/L7o�h�	6L��_�}͹��(!\����԰�&�P���Y�|;�9�F���l�%��h�5z�����Z:��j�B;U��cd`Y���|�)�x-�Z�"�2h{��:P&�sٯ*���28�O�q���Z�����x��_�n�����C�s�؝2%��d`\���6��� __����Q{{$v~t���=�?@A�0|F� ~*EQY����?LF���/��=�63����&�K.�Ȗ�_�S���0�'�ѧV��0����5��ڔ:��3�!��]������^���1pE^���H.�ݸJ������>����2�wzb��y��Ú4Wm��<��ku�1x�׺:�{{��F��#$���7hV�11��� ��2uk��6�ظ��+w�t����]ך&�L(������I��c�C��@ע;�ԉP|ľ8E���V}"L�e��g��%"����KJ^Lo1*a���L�J�v8qo���<�t��{�q�0n�m)M�.��9h���Z{+����� �sc���&P`���F��C� ���h>��'��{��˶u�aӱbyZM���)-��`r`A+����|*W$�:�$��&�v%��tm��y�"U�d���%��
��C����7ZL�rG~~?<gd����q�\/�u���m��˪9H��uj�Y=�����J,�9�c��ܔ�ϧ:H��o��E�s��Φ��Ǒ� �t�����}R�s<�W�6��t��a�kH�b5ܚv�3��A[b%3&9Zj.B����D�������t+�ev+R��1N?P*��e�UUܫU-`҈S���M����Ma�(�#��IHP�%vy(�w� �=�8��pp��|���{;.�6����3�Ᏽsl�b3-E�,e]ƺ{_�	'�1PO7�s���=��ga��M;Nvs�(��Wi��r>]�P���p1#���S�n<�31i�v�[�8�0���Y~����)q�Xfy{�O��`^��@��#��x�ws���C��~�,|�G~ҁ�mש39���]0��oAO L�*��7�˚�e�,gpl�ͷ���T�碮H��,W��e�\�S�S�7E�	�H�ǩ*"l���;[��x���GP������cY[B�op�z<T��h���x3�)s�f�K����+����n%�>�x@h����������(`����'�s�����p=	�����yh��{e=���9��﻾JR�v*��dr��[[,lr�ϲ*���U��ފ�U^.�z!�u�Aw�_�擉��:��sP�Pȁ�6`ʖ����H�K�˅��/���
=�D��~8���HsE+�]��΀&�1:��9	��Ad	��fT� l��D�I��8�N���L���K4��}V�x��z�x�?�f��_�g���e3��Z��,[�@�>�)K��"��"�9�f/V�(<+��)�6��"�X��PE{H�;2�=\n�A]@���ܮ�z�#{ʲ�o��Ðs�,�:��1�@c	f�T,�*xf�tq �x�lR��/����M��z�C���t�Lsi6�\�������4V����j�r2�)R��ֳ^K:�n�uD�m��V�E(d�G���%:� �x 0Ԩ�
6}E9'J��[3U7��/�^O�/���g؏ ��Ia�ʒȡ���(�,�.r�J.L�j�A|��a Kv��p����)���h6�,�t^��0_G�X	�����&|r!ؖ�Y��N�j'���e*S�P,��`t.�<Q$�[�yQ>�����T�"�^��mZ(j�{�K�5Ϥq$'l���B�4Nloۻ;�EW�UE�kdV�8�Ց�
��i`�b�F��C�p�v���� ��R����v�P����0�O<1��y��`�R�3�zY�&uQob��)ܬ	\k}��v%p�m��8o"�V�1�Dś'�C��{���k�{�p�����^���:�+�TW��������?
wb@�������y��f�]�ϸb�FZ�������Fu'i�%kKK(�B:��k7P�C��^���(�-ۿOZ\(ؑ�s�L���&C5�iF�S���'�ҹW4C$�C&�Uk�t������'�O�5�S|{o��#Hڟ�h�3�@��?� �~<b�ە�Z�����a�j\/ ���9{(�ӹ=���i�S�2|�s�������i��0�==$*��U�+;�>~r��3��ܳز�wq�?/�C9�"y�!@��I����M�d���c��K4v�7��t�m�pF����{��<Ƅ7Pm;��S��.)ZE�4�Nz����D��~F����<��yx��V��@�A�����6[ѩ��l�/]^8����okd6�`��t���D�eU�Jq��P2,&�Q�A���6+1Y	X���E��h�h]MSI�l��5��n�.}�֖ΐ�o86rd(iC'��|�N�O�F�Bpn�O��혋�:��TQ����Xg�?$�~�9HȞ��e�Fl6���y:��K<��g�g@݈׊������L���fA��ꂻUc��sn�;(�ͼ�s�+z��7Q� o۹��Tj"��&F\W��O��a��R12Z*����H�O[Bw��5��"v^����E��v2���!&�EA�]�;5qdS17�p����ϔfg`�D�9�Y�i�+�/������h!�S��r ���2eb�J�f��P*KD�a��m^.p�*����,eu�,���C'l��Ŧ��zS쁛��� ݨ4��h���&A"��V��&+
�8�(�n(��c��ق��g�a�"$��|f� �����_t�bS��]M:���@�XJ�jF
4�*���F6{�L�P�ۏ�#c��v=�]���@����rɷt��t%��� Ʉ��:��s�G�S-O�p�v���#�D��ESG��F��q�-��Ԛ@b~��H<�' 4Ƀ=�I .ņ���X��!	�#�D�pS�T1��\��%D�몕��m�kxN;�X��;�x�Ӓ^�8�!U�e5�~�����n�����~z&h�0eW���б�s�ml��Q�D1&P7�������270ǻ��`��5�Ǹ��"��=RW������@O�=�j�����p9���l� �~���z�V���(XQai��wuu����	Qh��Vbks7I��(�����%A�-�����͆��M�m-?ƒ%lWY���\��\�5�;�i�A�c��/	�/
&�:>7 ���ԢA�X�X�F�����Ŵ�<C����7�$�}�51����Oы�#�M�l�:VG2h�Up��#奖 G,q.ӟ
鱟f	���>m���5��*O�`��3�aS�䠫R�:�d4���R�2�%Y�L�`�x��ռ
�h��~0Yh[�A��ª
ڳ�^��s��4��|#�PIO���u����4�h����b0*�\ܿEkۯ}ޏ�}!U�՘�g>�����ɲG2��K�`s������*�m)w�ӮuD�1~�U��P��# ���@�U#9��x�?�����1i�:�ߎv�qR�^�'hp�5��p�׏�D��4%r�h>3��m��fJa���80,̨Z6���:�%����%�^��Q�����;��������
>	{�g X݅�uL��,���ҊSk=���ƶ'��8�b�����۵/�U�1y ���ы��wk�6���2��(x�� ��Zu�`֊.�P�s�FU��N�/����2o`�OU�v�1w�֫.���z+��Kٸc8��n�WA����z/4���ѠmR���u��כ0��,�����`�׽�-�s��)��X����]ܮ�ډL=ҹC�VJy&{��`����EuQ��c�bO��w���@F�a=D�U{ʃf�0���������%����gh�v\��[�.�Z���>�9dԉW`� o9���dܡ��8J �Q�i;-��b�������s[9$�#�<���4z���~�e��&_�@��K�(y� 2|Q�%�ᆢ�5*����fo�#}����ހ�����dP|�N���g�}~���zݏekEu��+���]8�xR���GԾT�W�]ٻ���"�#���M^�tu�	*�Y��!%�wX?�E9��%1�k9�SÛS�W>�,��c����2�%]6��a���L�#c�����RLl	�+{Ń�9?s�.yJ8s���Ď�`�B�4�$"��g�f����=�V�VF���]b#�����!��^��P�p�qH�l��~s~|�J.�K��/ő�o���S+�ҹS����~G����7T��Ŝ�U���I�|���o#+Į�K��[����uO�;�_{��y3_>����HTa;�&\�	
�����b���C�5�Cׁ��ý��!z��?�<Ѵ/A��BA+	��B�|��_�U�<K���)����7%tu�.�����j��)�f�>��۷�A)[J9�s����R�`� 
�T���x>ɸ�q�y#9;k��q3����cL%����u�h#*���}/TE�������ZB��Lv������8x{����H\oAȇ��1������;qnH��"�2B V���q�Н�7�P}K��S���}�]x���Raӈ)�7�e�Â}V�X���M�;o�e{�%�0~����Dc���8����g��n����ܔ����x&���,�p>�t���0]�v���m'���@k�n��F[���A���&�|i0`9�w����4ʲV��k���A*
��GJ�4�^FZ0��uf:Ե)��_�m9>��R��
a�Br��x"��u��V���f�ù̅I1.�a�3k�V2��	�=n��Y��Zߘ*w�[V{t������ʃ���s�羀�v���L�}�H�r�\��x�x�.T�e�Ɍ˗��OIs���eI�/�7�D2�fyn?���o����R��{�`�	�l�3ן�����o�1؈K�k����rt�P���d	�~/�*��B*v����A=4+	Wm�Y�����Q����'�y�_p�P������ ���#��;��b=���_%Ğ��Xx�1���2[��=)0$Æ֤縡�Ɓ��y��.^�M-�(����h���LdyW�0�y�6/�a��n������O�MOa^-���/��f%��7;��y,��m�&�fRX�d-�x�y��E8> ��&sf��>��r�%�3��3Hu���M��je{��ʹ�����S����5ߔk�Վ�3{�a��͉kx����%���ST�^�X�ʙ�*���0�v�tH�X�N���L��Q�����Il5k$�#a���$ ��?�:�L�|?�W�wgnw;o��#%J$㍦��u�fz;$�^�*ew���Vj:���E�n�ݻn2-�/��L�P�O�vk�(�L�"�8Ӥ��>�#��L���o$�������#;�'�z�HqH&N �}b�u��r�os��nae�k.5a�)ծ��A��Dŵ�`f��Fֿr1��ZA2�뱢'� Qg%��-^�0L�+ot���+u���+q�G|���1��.��C�I����BAp�V^v��M�3�D�6�M�ɻ�)�U�����j���G�m%մP�O����F��p����=��S�d����՟>Nל����D2|��ު���1�R?�݇@�5��|`�{Tt���P<ciח���1����3�3D��Cх/gΐe�
�"d[��L�|j/�E������ll��z
M� �F���� ���EVtLO٘�C��+;�HW/݊hJX,߇?O(����B暋)�|�������E����`a;�R*	e��Qh�C Q��E���I��O�gr���{�����c�J��}|Nt����o_�I�#y1�~f]<j�c��� ���O����[�%�l��8��$r� f���z\��T�?H0k���)1�C�b����i9�lb!����(�h�D�W�#�ʽuj�U8Y+	EkӸ�̒'x� 0iN*�h��M��]�Az{�_[�+xV
Ŵ�w���p�bA����d��}<>Q�7�%t��F��YM:���EwD>��ߣ_eeU�볜b^�Zf�CA� �!p���Q#1f��($ȈQ#��1[4���$i��$�����)��dQ�c�ª���[A�k˳Q�յӫ�J\����gϙ�1�;�|�H���Cn��`0�P�ր��+��=8e�����觟���Xw����'א/g�!
���1�P��#^�$
���v��cnZ��l���!2�a���\&t��@@W���I�Y x-���m�1:E�Zl[�/���:u�de�~�Xb4ND�g~�m��5��6EOc>~��Q�0[� m0;ن�e�ߍ��?�&&�G����F��|*�=XN�?<����=�[c��
=�1ec,:�!_��v�}>IQ�2/�cgf�~��t��G�yT:��Lꒅ9G5���f�I��a���v�)%�h���G����lB1wk�t�x`0�]킲���D
u��d�D��(m�H�n�:f�9��W���2""1d��#jhR�����ӿ۝��*c�
F��!�-(�Ӧ�	s�懶�)@P]���<!���=W����GQCw�I�r�[�K���4.�
�*pCMns������:���Q[=}��T��}��ϓyhe���+g"+\��>*V"�����!<�@���l�3 ,t>H���p �c+c��ۨ�#�݆ʳ=F���*׮]�fI�_�>v+�Ȝͮ<�z��=�
�	}���"a4D$p�ś��@ղuj7���j�H��(=�qXί���O�j�wQAe�U��aƫS�%n�Ґ=E�\�s<�hl�4@��af+Ё���f�o��#�L�M��k~%�������g��W�Ti�g����T��+n*.�v�S��V���_�<ڢ�ٖ�zr���o�������ujV�:1�%$��a��$yb\5@���gj����%��΄Kֻ�hP���"R4��+3�45�}.�:�t,DZ`�T�v_"g':�E�G��Oq�D�('GR�;�s�F��օ����v�!b���'�lk�b�����  �/Ւr�Wv\���NoB?�x�m�c�/xS1� 5����GT�&2Y,3�5�$=�RKI5w�:�"��a`rŖL>��#�Ē��8VA���>0�N�'i�"ӕ�Kca(1P"��❪�/-"�#}���):��>��f2�I��Pi�_.���� �63��fF��[o���%ͮ5E�N��9��:NN��Ú��==���v��v�����y^��j���oc�t�	�g]e&�"E=�R��#|��]�V��>�7㖀��fY�=��hPC3+��Ֆ@צ{�#םO��ӂ�2p�����ɼ�飑9%�3��h}#��R^���J��fY��'~�B���Hn���/�Y�͖ÿnꪊBn���ח����l��reI֍x=��_�a�iu$�0��W����P�[#����V��;��IXfs��B�X��F�<��.�Pr��(Pe9��LM&���q�e��Em�����?�VZ%�C�T��
�vܔ(/����85�_�	��W0+�E���B c���L��^7�dB�(N�mJe.�P�`i����/�	_�J���7�Td�NT�Y[��Oc 2x�I�ys8P���>V��xW w�VC�GaxԠ@M��b��"��p�]A���{Gr���Yԗ4�ޏ,������Q���+�T>�1{/�a^���PY���p��bVm��E�0�d1nV;(g���h���nnΈ̆]���To���5�CP/w8W��F'eIDΥY��F=��
uɴ�aTO
�F�A�h�-�Zf���<�BT��0�^�ǚ9�B�3��+$��ޚ��1����������1B+S_�v��2�M�W;!bɤ#�P�|���
ǉ�G����y�S=�y�~�j6X�p%(�ˇ]a`@~2������1��ڧҬ���r=��[$m%�
�x=#gٰ�@�SG�2O��"Q�&L&��0m���#�S��Jn�~�i|���[OO�t�cT�/�	�܉Tpm�[-�=m�0ѝ����{6�(=��JEU3�rH�V�h&�_��*v�?��}?��2੶r0���LD��+r�>������+p�'%;�ńö��V+�L�^#���c-�ʩ A�W�*��ɿ�6Ub��>���.�aK�(�jOי��$G1
 p^|m��]H��IN�%�CП�����w�����@"�ڲ�)_�[W�@|��ə�d�>���j�����\���#�V�~�/�
S.4)^�AGN�����_��3@鋌�@/�)�l� �ci�RP�B��jZF�Xۥ�x��o&p�P
�t���iԌL��j���*au��,%���$x��C�v���k��j�0��+PpKULx������葴���_�`(M��nsB٨T��y.TV0p��U��)��C�gb����c������0�00{u���������f#<{��Pr����%� �`��{?X�������.Gܯ}����&G���_=����qY����ãt��H�֠��rI�-�s�QZt3V[�$��{�ƷJ�Z����?�����D#(Q����׬�)��c
� ���$�g�NO��1=��qDr)l��B�i�Ph.5Q�|�G��Y�p�e@�1"G� `�4�T��qv�������W
]mm�\��Բ_���1wlC��!�����B=����s��vU^�/�#���G!u��`i����Z����P��
9R6�:Df�����-�8ю�Sє�*~$k�e�
��r��VND���P;ɻ��-��М�d�7(����j���g>����o��uZ\�.�׏�MM�quM0���2]�5ǯ{E�5�{<��*�v� c5,LfT��� �k^�h���=�B�0�9uM� j�e����ńs�{{�EŬ�����K3aͲO�����~�s7�nܢ����\���<��;ˤzII���e�\4ɧK]@+����-L��-^*~s��r`�q5m`:�4^�#��ցhk�o;�q��{�v��K�]�=�2D9ʲ�T��m�N���J�CN�����.Q?C��ٝ,�E &T�*;�	�f�]Z(a�a�#k�l�>#Y�B���{���-�~�9�U����>sW$��^�yƗp���5dG4�Xۦ���u+���w�i�������	fG�����s�踻�ٍ#��A�5�W�=�~��}`��l�3;��X��a��l�~=�@���v7�z���·|G,�V���=d3��sf���F_I�|�9�ͥ�{�d�?6�[�^�dGӵ���GrM�H�o���Z�([(E���թG���f���P�Q>A��W�L��:.��M�Q���,%~����x�܎�O7([f����ޟq�|������u>Zݨ��x{�t���j��~�����d"�?94�iy��:x�/У;\1T�z,��݆:֬��[gݓ7�eg	R����Y�$�͇�c��׷ɇ�G�a��N#!�|�q��P�XPy~�Z^�L�,~��z�٪W��R�\��ȫ�o���pEz�̍:�V�
11���`%n��}~�f�^��%�[U0HN����Z7��p�:��߽��m����B�d�~��。s�6l�� !<f�1���w�|VoZ�+e:�{��X����R��8�-/Y��f��z���t`���E0�Xtc�W�W>��L��9�4�H�:�v-H$��)�XR[(�)���v(�<����} p�"t|�	K��}�� ��wN;3K���Y��u���s��l�bpI�|�������B���Y^k��a������w�/��� �¥x*$JNN��6PsP޷���k���u��E3����M/I���~���yո�dT ���N�ߗ��
����EK�E�=��ĳ1LBo��*rkJ�`������@r�_g�T�����!��6ڹ���qk1WL�Ȟ3k�jY�9��@��_��Z�\�CY�	����ச�`\{�y�p�kj�܏��y�9�C����s��Z�wa��lv45� K���Yr|��x�����
;��O��<��ԥ�vAo/ف6��~��U�^��qKŬ`��A�r���(/F)Sw�N����fǑ2O��b��� )��1�f7���`�'��q'Z��ɤ�]�chYF�XT��&�e3��)M-���w C�)6�h��ڔd�qe�����O8��0vewk���d��s�A�����ruk"��m��T�֐���uיf��危S7��� _����Z�NR�35�>���^sZ>d��!����P$.2չ[/�f�g��J�v�d�Y)�\���\�_����zk����}�ѓՃ44���߄_>���F�YD�⒉_m�	�]�a𬩈���%;�V�����z�D[�f�j�����t�)�J��M=�T$xX�D�H?@�"L�]�41��Heѵo����4�c��� a0���r�h���G$������0�̨��3�TߒD����.��j١�0�RԦo��G]ů�x�s��u�/ӈx'�ԗ�6&V�)Ȧ���U|k"����>� @6����c�nQ[E����1_� c-r�u��,ƒ0�^�;���K$�����e��+o�q� _����NE����9����%�=�C�������U5�W��)�l
��5	i��/u�S)߶P@e\c��!�b�p޽��Y��[Z�Ȩ�h�\슃�D.��{�"`7j4ai�»qo<�WS�����[*��;�b�T�U1����|{�m! �G�2�nW��cOmJ�k��'�Ծ��ַ��ғ��i�CF?���m�
��������$���#�YJv=�-1F��[<�"��CX���,9i���{�F�n��{"M��N�Ff�;H	����t2�_��r���8��檜|#���M)!������|�5z��tí���Z9�d7^���Ϻ�bD�y��CRj��]�G2�3�K��]�W��V�r��h�:n��~q3��+c�
��BؤQ�E�U��i4�k��w��R��^�W��cS�{.�&�O��$��ظ��E�����"�~�4�j��|H͔�M�<�h4Զc����v�ي��?��'��C���cf�N�D�-�e�
��ǁ�'6.N�����B�	�g&����O��D�wƟ������Cm�5=��ߑ13|HXv[q��
I��Y��u�x�|�~���T5h����Q�&�^V~�j5�\����w���.bf�{�FSO��T���{�R�ɞZLG8�'���0�Do�bC�����m-�g�y+��ϯ�/s���;D<:��y�ET�~�GI��l�3%޲�m �7S3�d܇.n �Z[�!b�[AL��-g�J��^f�$��m�i��!���{ը��c�5Ie��dN����	�I�Ӽl�9u"�4`�5�r��FG���:��2�����Q����PQuR]�eY�j��m���"	q�2lB�>d����e�U	��@�lE��	�4�vl��0N:�b�+T�V����ㄦib��ݬ�\�>�М0��J�9��7���r�-4"wxir`�i�~���\�ԩ���s�L�������M��/MB>K{���hR�$Ԯ��n-kó�ww�z���b�+Ү7�¤��&Z�wu����ɑW��ĎT�T^���UiK��?�rȁ�+�� y�UT��م���fAzt`���sN�7=����t�I���'�~wYp�H!��01�S[��>nb�m���T!�|H3�1J���$'���i����@�Rm3��Jߒ}���n�p����؆�Z�u��X/�h&J�#���FS��մ��KQ�GA��dB�e|�u��y���&������r4�%Ħnm`�͌�K�l��;+��T?�c�E"R����&{�nC�&^�]TF��6�`j�1�l����hs���*Y�,~
N��ȓ���QmBE#��3�Z�9�)�7<u�v�#Qд?j���̏��V�edbP�wZlȩ9��$����p�^PQ�'�����΢��ضylj�i�|+�n�pm�㎒��2C��Y ��-.v'* �ϴ���������3Q�W�z�Y�T,a�<�z+B���̣n$���l���1Ӹd�!���K��r��FS�2�0\�:�"9d|�����J�����F� �2$��!�d]���K.���9���Z�b`����e6��7�MhۆĪ� qFr��E!kg ��kK�q�js)9t�eqGJ�Re�8����`V�d��
�5�E���O�Mi9��W�A�	ۖ��A�����'){f_J�>�>��c�y1�fV�Y�q��N:2����W�KO(	�)OwFt^@�Y�����[B
T{��D���哛}�+�1����,mX׸�5�%$+Z6���x%���T�9�g�#K�����tC�UH&:w��º���T��~��W�R��H��z�i�7/O�bL��*Kq$�dt^�q#e�U:_<Av�O�^�"��)*�҆j����ݒl���@��ȧ/2�`t��y�-�920O��-��@�?I��-��W���b�����Zj���4A^��!�<岣�s��f�̯���E$f�q�̦� =���|�U*�~I��K�'��!Ġ���,��V�X�xهò%�ͱl����F�KKW�Ӓ+���(��buנ}A�[R;��p8Ͳ)8�&����hZ����Lv7fP�M����������V	�E�m�dO�m�dM��d۶�l���n�d�:5Y��������/�g�k����o�}7�<����Q*&Dٵ&J$ݴ��SL�!�0Gi���z?��4�3�r��2�Y-�� ���j[�r�z���;��L�8Q9C{���-���$��AF_�j�Gz�$l%|ط�+=8�p�Dǁ�[(�Q�)���_JS��z�q�����\56?�����VV|:����9݌�`�7�aV��O���M�"0�*�nO�0���Ј�3c���imVtvǗ@F� i	�=���Dji,X�Xa~�e�4����*�9�񶭶lH�`��z���du�Ҕ^�Y���Se%;B�-����\VV|)�n��/n5Yy������b�V�J��� d��o�F��h�:y��$

Z���9 �6�����b3���1_���VӹB��_�۽i�(�Nh�f*N�o�O>d�+�1��J�j�憓���[��GDq������ga���E� M2$��d��=A�Ư��;�n�hݰ_�9� ��\�~'Z2+��t#���H:ٮY��������=w��Ŏ+6�؟� ����/��ML���c�[k~JW��_z�]sX*��]Y`�ƅ�>I,�@o$Bc%�#��@�&$�l�M>��	��ZR����;�c*�HX�3C�O�|��S���,E�밖�	PM�T��ݳ�Ű8�r&X���S��n�ѻ��/KZ�]�i�]MU��$�Pzи�����Ca�A�}�BMi&&��H�2Yf��:�?h���v������ӼD�5�AD0r�rA.!ά�;��b�p��w��ڂ&�B�(��@e����k�,6���������e4~_�X��h��g�u�;�3(��k�:�R紹k��p)G�ų����/#P����t^��)��
��N��`��0<������#����Lo�l�I��lr�"[��M��v�$�=�o�/��&��v��6N������ę6��b.>���h���)&9�ܙ׺�������i˷��5��Ґ �fLޑi�`�q����ɂ�[�s�􉇄d�0 A�(#��b��M�^��t������TC�I�H��Z? B��-�V{C������k�-�bV)�1չ� ��-��!��k
s4��c7˰7v�Նv��q �������e:44��p0�X���j�cl\��Ƞ���GY�R�8����1n�ޭ]}x�������;�>s�;?�#y��Ep��$����F��Y�f��o��g�1Z��ct�UN5�=����\�ʆ/�(���'́�6��d�#�cCs<J�N+	�V���:P�/���02Ҩ��]H�^�O�߄n�_�;�z�{�C�������-+M�3	n�և�ǿ�jѾ3�����J\����G�y���]^Ws/����wj���R���� 6�0:{�c���gĲ��p@��!C�Xy]w{y����
��/��Ӧ��+��x�Ŗ-=m{WL|l���޴����^G����|������{I����݊�
�A��؇����Η����ޜ{��45 n�}!��E��� .�rn�1�rZ �?���֙�~�����u'*��>�ڑ�^����պ������q�'����Z��n���0x��F�aa���y�y��0>��3�sf��!<�M����q4G�/�X�=�]�&}�ؐ�,�@b�t	��d���k��.�B�1�l�d���F���|��m�@����c��~(��y�Qx���O��W��I��Ŷ�����+��vls�p��U�9��[ե�0t��@�|��+Y늙3���� M5��F����o��ss�Z��Y����Tml9+�~[�ܚ��ܮ��r���a�U��@�k3�h�~��H@��O�Ĺ���&��|j)��	��-,���n���P"x���D�Tn����H��r��7�%߽EO}3��f]D,K'
���'~`�.c?2K !K�#���=��%���:�i�����c���3���1KB��Y�po���u�F��!{���1�3)c��P�W���A��?���N�>S�&41�"��|����;w��M�XV�Y��i0��������n,��@�JkH�w�Z�;1��r�zR��2z-Nm���x������yj��Gu�H�VUL͚ɠ��~iW9-��F��ފ��Y}s����h�����p�Pң�ײKO|��0\@hTv[��w����5�^����!�s�����c���d}����a�u��=)p�뵬����
�K��Y2o�!O��"���|��7ע�h�V�z�x2�����"�&X�</��T�:��q�*�-qʹ�Y�ʅ��%���c�|Hh�,��в������ן�Sx	dCrl��gY.�5�2]sw:"^�	��1O���6:���+}O=`�y�G"��j0U*�����Fj�M|��6�߰s]��u�F\]�>�c�t� Vx���N��R�ƭi��@�����'�a�-��6U� T�)i�r%�%�~�6D��j�ǯ�F�EWBC�5���W�o�ˈ���ׇͧ,�C�B�l%�눋��!	���E���x��}��yKO����$y2%�K���w�c��J�}���:�Y$���	;�Pg�Om`,$J\�4.�on?|�T0G^����)[v� �F%oEz	�l�#"��g5�!� Z��ߐ(Gps�ke���A��f����s`j�!R��=�C�Y�f,�����'"�4�Dnd�z��5�nR[Y���0$�c/�Ն����O�̎F�Vs����~8�i�M�v�l��"q�5����Ie��i":��͔�J����c|��IM[]�5��u��oMu�+(����]�ev�\��t��C��M X]�؋k�\��MA��%��v@C�ͮkW>�In��MJi#N�frϑ}_0����\�&Dя.��͗]a���q~�/6Ex�|c�>ʙ�\s�*`����_��`�*_����E�d�H<x�5 ����?��i��q�n��8�V�?��'~��Md|Y�c ��̴.]
g�gRN�?��Q�d�I����^�������ZHr��0�HEb�f6$�4�X�L�M!�+#4�>����DÓ��]��)z]*w�w���8�<�&���~��{�:�0�$��G��ҧ�S��	�o+\�I�HTb������pӽ�[5q\`γ���zb��Ń��ϰ��z�ţ�>� _:�����*�sy�n��ñJ���o�2�<��H�=��g`�[:OSSRƷ	<��DDoHZ�+Ë�xqh�l}2����H���H5�v��+���_�e�o~x��J@�9Q:Ziٺbn���r�?I�l.�e^��9���d��ި�뉅�����W�Ѽ�o��4(�cL�e)����CQKv(��:z,YFL�Xj'�6\ۉE�6>y^x�7,�_2e�t����KZ���R^�|���{M���ިT0f��J��:�O�^B��������?�O�'p�]�J�ۑ�G��0�^�U�Ο&~x�3����D���_�l�І�J�FV�!�Qe��^����&�IJ��L�6</U�����lw����*�0�\�(X}�w��~ש�����ǞG_D�9H��g�0�
1�o)r���s��.c	?(k3�!��6!����5�,�\�j�z~��tjU�$�)������ڟ��y�^3d"���W���Gh�B��̠d���"��(j+4��c)�&b=���=��w^��Z-%c���y|/���g&�Wϻ�����[}�B��x��������+��/\�7��S#$
M���c8������*��Iqd=�xB^33llB��:���{��wPJj�HXe"�7k}��*��@5�S���c����!>�Q]dA>����I�B���N_�-P�";l�P�eH�TK��X���hg���;��p�}��4Hak��2!�������mzy#�0��.�BY[^6�o)��Tt�����SEx*�?���@�?%~��sK ��"����,Yb��ӓ̜Q�ê�������&�l��@-x�6����wr۸tbp��Ի��Hm��9���]|$�
���bS-Ap���h��I��R��=m��:��l����~�^��f���),�w�O;>���J��Rϸ��~��	�(���S/~��J�$��i�Q,�q��7����*�~�/^f*I"<�*�D�t��'�L����3�`��&�z��w���*�+���Z!�i�"��ߴ�Jv���r%���0���/^�| �z���2�:��Y^l���W��IW�jit2�X�����N���77�KE�����F�z�� �'U�
%���kz\�4��V��xu��l���g�v	�`r�נ��db �hHHL�����L����=o�#�<��?Vw*���{�D�������|��%b��\�T��=�i��%��"����Y��Y�����|��i� �?�2�t&���=�<�2M�o��Y|�ގ4÷��ߔO�%C�2�M41:A^5a�m{�#���W.;�e�"JX�Q�b��؀R�B^�1u~_��+2P��gF�x�P��LM�����(�X�C:����M
���&ȇd�gU"�/�n��*����q��m뗷���ɤK�CKQz�Z�nv0.��N��KX��;�ZEz�J%�K�l�O۷W8�;���y��B�j�|��%*�SM���5o��9���X,��c؝'��x�ymQ��n3�ӊ�`�1�4h�
=Œ�\����7�� J�r%�]0�#8 %�:)ܜ����=�א4aY�V�8i��Tq}gߌH-E���<��d{�;�9s���Z���~>a��>��g����k�	���J<�i���^� D��v��6dK[gԗ�cJ������5�	]>��5t$4�rn� ��O�<��h��>�q�h[�T��$��������I�$���M(<��Е�I-7��Ĵ��؈)����V���u8��bFD�݇$eX���3�j ��������ŏ4��xyy�M��.��c����Q���%��q+#ہ�2Μ��� ����lM��"݊�"��$���ݛcN�����9���	�y�L��Q��.O[2|I��RU=ͬ)Y��MJ7^Nҡ��yw/�J��4�Y���s1_��%�ȶ"�>��*2̼�辌��j��T4m�!4�
��O|j
��8�yJe��z]
��[g�ny�e��YK:V�-0o����r�
�u�ôS�O;[��U��w�a��7��p�q;P[�h9��cH�~)d�ώ@��	�⁢2P�W�u���?�c�j�u/�g�	�Kvi0,9��5�� I��xy�7 4N�Adj�b�{\s�i��Kp��?*Ys%���gr�ʗ�d �ꘋ�@SԈ/�������"�7<�>�tu_W"��aC��~�O�f0��G�x�>�/e482���W���zR%sR1����!��:�1��H7h�+-�]��1�j�W̒�K��G�4*�h;Ւ���m�ץ�E��.���態v�˙Ҹ�0�`�����l�N�MzT�I}i�z��0�\��m�#��b�yc:���@��u�U�f���P��7$((N5���ע����lR\lTyN��Iz��I�1��Z=��,���Zl�7�6�Du�;ol�E��9�̷�%J��o�>2p�P�\h��ژ����C\�[���M�v��G�_c@
�u��,+��X���D�料K��,ӹ$	3\�&J�`
�[h�Y�娜�a�p�t'f��u�4�^�]-��T=�z�$���ѹ�OlJ������z5o��)P��x���_֬�钮��G3�6hGVƮ�̈a����������z-���R����,8��������'l�5I˻��	ߒ�ˡ��r�`R���@�3,fyiɧ��܁*�mP�"u��H��}����-x�/Exah|�=I��!Mo����ml���� ϖG&�؛��N�ޗ����� FVU&K|@7 ��t��n$���rd�D��56ɨ�����~�J�n����Y��R���Vgq�+WS[�t:�
�&z�֬L_�	��$�{3��?�jaQV7�B���D�g�̾�
϶I	7��ѐ��g�Y�'��o�>?W�3Y�f��-34��`p�[����S����RK��yi���e�A����ȕ��mD�������?����'#**x�@޲�� ]�_9�_{��6��<�tzP�?OO{�8M�Q�%���P4�z��4�ZS����	*=�pY	~iVb�n�4j�pʍ.��%�"��.�zTD����>�	�¾j�=�1�-Q��s��S�]�<�a��E4XN�!{��h�Dk�#"��7�_��ĺ���Q���hbĺ�WCb�Ŵ��ۋ�b%폭<��Y�j^�3��0Թ�s]�r�h]ҴU�ϠsW9Z�UW�_�J���"oZ�x���#|�do)n6֋�X�LCx������G�3�EeXN�=�D�����7"k���Ai��%Zt^��>4����n���Re=}*\]��(��Py	�^�ը�e��&m�-�ʎ1̥$�����N |������u���1A��3�6B�c�^ots�#�4/��uE�$�~&O�L(hE�Mqh�@��~f�B�K���Q��/~d�_�"��&��_Q���ԒyL˛W}Gbo�����<Q�o\h���c����{&��K�Q���"p�d{/\r?�u 6�v�#�O{�s�^}'���W�U��,w\�����֟�������^�e�z��?N
�zW����nM-�~^��?��r]��I׫c�.	O]W�W7���ge�@��%����?�w���h�|X5����d�dŤ~��V7b�po��<w���Y�)��QA�)���A.R�Xn�;��m��-;6m(��{e�s��"T�bD�Y�8 ��Y �y��H��ue؎��=-M�Z�_��g����*�2��>f'�ۦdg���\�����6jf���i�"�G���ʀ��a��tI~��S�X�|��뮐���H�'������}I.�Pc��l@2��{V֕"x14(F������^����|��C��,R�
�_L^��E����w;X���g���r�5��S;w�A�Imx��ΐ�ï�2׽�?�T%p�[@�0\�9���rpO�n�����W7���i���}��1i��6�h�4�׾k"���Y��`;��
�!�{�׭D���.��_Z3wi��8f��b���X~�Qbv$!��.��!�jZ������N~M���*�׆����[����629�G( ���!h�4���\�G�y���9��=LM�f(`�r��~3i2Ȥ���s�A�8�8{a̙�<[��32^F���V��o��~��/E���l?a��m��w�Jӆ���<�4�l�}����ˎm��y7'���|m�M�y������:c���"��1��Sym޾����D=�f������ݜ�e��	g�i��6i2�/�������ƹ�ވ>���*���4	�zPr�
V斓�F:!��nQ�Y����}q���!(A
��0`S!ɴ�������P�U�h�m��4�tk���O���T���m�9�O^�?쌡Q�H�V��B�3��f��:n��}a����z���<8��1�?=���W�?+��kr~6���������S���i���Hя>��=�z?�:��k���©�@cwm����t���p����
0���jA��":���G��^�����^r����s��������l_t��'�+#�d cC�:�V��+̝�g��������(� �<ɍ�{��Y��[�;q�xN��0��J6J-F������\y�B}\�|>jS[���7�������O������������.gj����G�_I~$G:�7��Q�Y������'�Z��kP��W����Q�n�zm�����"ev0��+u'�=JgOv&�2�IY��բ�63B��|��^/]u��"�+6"�A���r�:�X�E��鳭~ ��3k����z��r�~.�I�����1�`�y�t����-��4�~�%?ً�(�l�y�"��&ͥ͸�3�װo�4�i���HYپ��$�ж�A|���C�]]wW����
}�1O��:/u�G���is
� �x�8!0��E���iۃ<spZu7��:�.�"�x�@���U�_z���L���Ev ��k��ȓ��ѓHT�{dҗ�k]@�qO�	��6�N�	y�o��z��"��e�����5�YtJ0,��������N�R�]���sfx���F��\�o�\DQ#�U��h�"�t�~�3}�ArURgn�?��JrDS�����{��rț�`8�J9�+�@^�9tzn[��u���G150w���j��M�W1���iV�!��8u,���~_P�Z"�A�2EՈZ���b�C�$�R/��h��ܮFg�Oj3Ә�nz�0��0Ҽi�XM�� d¹ᒼ�"Q�L �����Kڐ���s�,|�@qi�K�qGWȃ�a5�!�w�����/���=iE�s'���В`�:�?���5q�|��83y�GEs�o�R�\��Ȩ}��� j�5�{�J��:�:�q+J�"0���ct�\s�ϐ F��p��=����k�,D�M?<aC��1����kc���k�$Z�;[Xa~��"$M��V��<
�gT~��w����	iO��^���sN�Rn}�tf1�"�%
G�ÎVZ�cr�O��m��9�����>?z\l���
9|�HPpK������Rj�P ?��(E.��h5h��0��0�1�1��Y�x0�}Xԛ��x��p��6�L.�g�mqR+���~�)�C6�����[W{�$֦A'��#�2��lܮH��ף��K+f!�	9�A������b�E�B��Ċ�Q�3s�>.�L��΄�F�J�s�j�B����0�� r�pÈ�5�y��k��5X�4m�	��� �-�ٟ�Qm�٤^�܍Lk�. �w���z��Z�˚���1�X��u!�aӡ��x �O'� q�(Wv�p	0=˫��^^B�����L�q�фB�&��V�0���w<�2�"fm	#��^'W�dYy��NW�?M�R-�/شu��$/�hK�&l()T�[�E���aשְ$�T���T0�C�ǝX�f[(t�� 'q9LE�n�����ͩ���J|v��Z{��+?v�\ �F�Gx�	>#'|n�Ӓ���Q/	��FV\?3�RY�	�����{�M(����[(nj]�v��!�\�/���"Z�
��ufF��^g�	��J�(F�G�p�E��I����#8�����SG��fx����!�Ҳ����"�4�2�����C�� �N'V����V\z�quX�8����tP�f5��^4��$W��� �.?���f���U���N���/���u�� �=B�=�]e��vE<9&�J/:DEG\E"�����?j)���.��^���EWޠ�ģ�,!��#��׮��i��"���"*R��������R�c�3�����jU5�ߺ�'��� E#��#a���J^o�����䨑`(	(�r��KjE�gZ��=��bV�q̎;�<�N�#ߘ�<�1���\m���A��H+��:��B���v����hZ�`��`��c�
p��U-�"E��� G�K�cݟ")�dRh����a�,�Ȓ��eĠLarL�C%��1�W�����y(�E�s�!Dy�!C��a�K��'��1��q�i��:]� �cUn�q�މ�l4?4���#X��4���5���F�2���k�I�,�}�>�·��9�22U��$i��GzD��Z,�=�1�!u���$s�9:�8�ɴ<2wk�6A~�.���g����]��h-�(��L%R�l�6xwɲ|�m��� ��}��)j���t�_jf��:��iB���������Jza	-�8:-����Ky��j����G,.A��JQ�2-p���2�<��@u���%� ;z]�H�_AL3�a�����o$���V�/��d��*�P�������2鼌g�F�'�:��^�/���^���e[2�҃v.n�K^����|��p���\lAXL����k�R�v�� &�F�4Ȑ�X~�f�̫"uH����_Y(�L�������$�?t*�BԞr�6IO}�/����uz'�*��_���R�Q�o��8�����ӪM���uM}R���~��qŐ*�S�?�����f�E�����.�m8T��O|*��OK2E�zz��ǆ��Y�5�:.��E�Q���ˬM<H~H��VҰ0}������-�J%Ag)��=W�2��{�O�~Z�����%���֙噏�2���Cɾ��]V>��� ��w{-�LDD��
�3�7[[�Ps�skE�I`W�/0N�1��xZ�n��%��q)��/a-�Q��[�D��OPGm����jO�A�G�e/�6���'��U�n�f$�#��b���AOr��G�s�Sj�s�L'���Hf���� K�g�K�>jX6�\;ZVX	W��y��������֮
��	5z>6�@@&Lz%{��M�PD����U6�]��Dh�8���VA�4��HE�ji���[��u��8KG�yJK�̤K5���[A^����#�EҸ]�l���H2�e�F�U���e�{\�%�� ��M���1#�Dĺ�"ܵ�Oq�G����X_K�{��`�7�T5���������y�4Fr��Y������ā7�g$"3����?ߌ��5�C�e�u��?�U(�F�Mo�>�@�M��&iۚ��ȑ��V�K�l��V�cF�h��eG�������\���<*#��8�s��C��7�N�
AK)H��у���U�U��λ�@�9�<E�8vD:[����%w�H$Z���<�Z�|5��F����,��R`�L֙��Jso[HZ�%�0�Z�D��������7�6��b |d$�`_ԟ7�_?�
'�X�&�f""�fWV*{@�zr,��Ӫ����?�؂$#ъ4��'G��Gɴ�6̼�ʣҩ�j߲ �����w����3ӯ�ޞLY�n�Qu����]Ĩ�|@:,�h�����F�]7'%�LE$ y_���j�45���.�i�0S�!(�e���j.�R-��w9"��n�����vY����&[z��N��4���0�~!������" ����` �f���G�ql�`�
j�`����?\ ���~y`���Ъ=���h��m~�1$[�B���V��ss��c��"�����RƝI�:F�V�;���g�xj�82#oo8MA3���=UO��S����5��"�&v�3Cڅ�1)K���f�K_�2;*�M����:{�+j�AS�a��̺�Ƌ�G#�.NBxu�V�u[��������w_��b}KԌ�9&!nn�:E)��.o@p��Â�Up�A�yV�1���:Z�-U2�.�b1��G���=`(��3�GD�k���#�5�XFh��´���� *k�?6����v1p��#����yJvI��1���Ĕ�\��F�2��$�t�L��n(�SL;�8A3;>d����GG�,_Ҭj(GY���c����G��"��L��2Y��q�):`7xu	��a�M�L�ߩ��-�KW)�f~WFz���L��2N��&���������?�DfL���K�*`NkibF��t��a����#��*��+�h���-�����0�[�׿K�e�7h��
�U,�0oI�G�8��Ү�wԜK�dN��e��!vd�_#L[�Q�{xz�k���ۨ�?a�K�4���E0[6����VUY9�`�2g~[P�U�6��� o
������j�*�� y��1�mf�jb(��/ɕW�ZJV�V�ڡ~.IZ��|}3Y�-
�cݠ����,���Q�t���3��{os3�P�3�V�D�v�s�]c�%MX�.��%G|��y^Ɖ��6��ԡnT��`)3����*>���:�ԋ�*M{����[&?n;�>�������3��F:t�2x�����"���2�_�ő4mUc�%�]��G�&G�f읮��ֹ���z�٘��'����á�B1X��rZ��]�F~9�!8:��p�=�Aߍ\�L�J���7�˕;@[�P�v�5�Y���:|H���gg��l�����Ź�۩�_ ����	;M
�I|�P���O��
~�\��W�?�[[WW7-��j�֬&��&&qh�z��CRWM�Z7�ot@|�6��5�ҼJ:C���XF�跍�1�s�O���nE~��q �Ar�/�[�~����������$Eq���3{��z\�.�tڗ�tP$��^+��9J9B�r�$��� Q����0�Ći�|�,Ί��#o&���@�7�
��N�40�%L� xX�֔�}�&S31�''͜��S�\pn�ABS��CC�T�!VM�ͭd�}a7$
�ͅG?���n��~k�u�"��yB>��E}�����8`�S�r��A�������`� ���N��-36��Ɵt�\���_�ו@���(��e�7nx-�������7t��t�֡�m�S�H�vJ�x�a���𬿆�i�-xD�+�W�2%�{�0�0k��O�+��"\�����P��@=ZH�`p��:j�΀O�*JӜӦ���������-��tqp���9��&�ۨQŇe�*��f2F�ME�[����܅�y��w��0%	��j���F�������Kw�>pq6$yy���R��#Dʦ3C�/�cx(�<�+[��t�b��F��b��Ъ��K�RY�b��l�1���wUӕ�^�	j�q�hm�����P�3Qk�ު��;��p���I0�W{�]�bj鍊~�$uF?�k��ڶ��R�	�������9��P��$�����ϼ|�\qLر�-N��b��_X��-S�}��Ok�;�#�c�3�����4�4̿T]8��8���H��v86�{�3��U��KF�Sɫd�F�cUqZ����_�B�r�py�E�Ey��]���Q��Q0Ե*H;�$l��"b�ϥԵ(
BG(��'��,�)�\��$���Q�WH���@�����f�.7�C������\�+�v�wdH����&�Mp�cLon'�̝�B3�=�j)�	�e���>��ۘ��Ybs �2��V�*� ��ǩ?R	S�����l���v�I9���QA &�c��5����S�C�f
6E2 ex%�G�x��]����r�_���dBSwj�-|]\Y����T%���d�S�+Eyn݃H�Y���K:��z�x�VMm��Dlt����|�ơ ��Z�QN�����8��?,��[~����iV�9M$Wi:}�Z�>�Rϓ�JK���ڕ�M�֛��{�(�{���!�l ����(N�<$��7�0�[j�)�T&�n�����bOd��h�^�&'�Ǹ0[(AIX�/0_������qy���bMF9�m��*�!�0s�w��\�λNP��"&ɨ��������:�E�aY�\��j;%�v�/\����E�d��%�0N����#+(�E0Q���K`�ݰ�<'wt(#/����0"�Tv�w�8`Sj����e��.ImR�jYzؗaD��f�(��)j�M9~�ԥVH�²֣�a�b��t�/f�l��8.;�E�6�����қ(��O�+z�o_����D��Ӊ��&�t��E:���n�1���ƺ���7l	��X�0�doJ�o��٦o��RVI��P�,����ڄ�^�4Bd�pu���Y^��n��̽25�i̪�!U�W+���_)��C��pc��r5nX�l���n����LX_�]�i�C���ű�=�H8	P�rY��'��ٟ��^��Yb�93@8+�,��I�P�I��X��)K�9��Nn���ZT�0��L�dg�o� ������v�����<�<��� ,��k!�,GCLADR�j"_��z��ozؼ�x�䥣�n�=���_��u[�p�p'���|�$D��z�Msg��dW׶tG���3{cm�ِC+Wz�ng�J$�P�	�)r��5�hR�����.��D�p�?����+����W�����~�u��&"bs=Â9�i�v��`4$=����:�z��8��n�$�~�+�ba���4C�j�WE�M��`�K��	s��鵘�3�t�����-7�Pз�Y��Z����U�A1�F8�W�R��N����z��9+h�Å��8����1�tI7�V��ok���'NV�G{)�?�mxFQ �L떝8�7�NU3��-j������`�+`�|��p�Z!�Fw$:�sQ�׸�!�-T�߂��ҫ��S;:�N�d;��t�$(1|u ���l�Ӵ�&�7D�)B�^�nx,v��؊���1��D/Q�*�g�6`�D��es���)�ш�(����F@��"���.$���Ȼ1O=d���$l�a�O���hN�i�{�.�Y$�oEvYk��s�����6�ls����½��-��<��Dt`�	��ɨ��p�H�at���NM��n���2�##��X�������O�;(�I�q��H��`�2[(8�P��'o&
�e,V�@�Ł��2t�Bs�P�	�\�<�+4V�f��֨%[�m����nRu��b��t6�{��Gk~���/���>���4���$b���zX��7��f3ǿ�i#�*vot���c���R�.-�x�:u�D3�R�>�3�����T,|�0��� O%"ȓ����e�`<='/�<鐤	�]T-Sr����aŕ��͐ٔ����r�Tks���WbM�j���m�rlr�)�Y��i���'�KתpSZ����'{/���¬ohgq��$��P�^#j�pH��K��Հ�V��,n�~��#�k�O�� ���4�{OOd�?g��ʬ�U��y��r�t� e!
)AE��
ƛm{�?l�M���=RhY����+�D]_q� ��������"�K̤.E��lO�wLF��҆n�*tj<\���S:����~�R�Xp�����ÿ�gL��GFo��ra��l�'���\��s�ΘRFSW�"��{�c3��<����?��M��V�z>�P�l�å8���G�Y1){�p���r,�A	݈�U�d߬�T�~�5�&�&Ó�Gu��뜱O"8���O�R��Ca�Y�<{�^��Յ-����k�"wS�����������#�n�ď�;���b�9��g$
S���(��Sl�~�
W���I�x�A#;�I�0����=��#�����6�/&��ɖb�����wGHK 8ט���~2������uRJ�b6�ͩ�&(a,P��8�l�+�%`=��,"o�
Q������\�%O�?_}���ފ7����_�����z���l�O�P~��f&��x\P2ޕ�L6M��w��8�A�:���0x��x�����Lk���~�%���3*���,�N,Gm��?��3�����I�n��)���E�6���]MɄ�u
�����̇V�F~��0;��T�0D�e`b�]kl#���e���˾�qp��ks)>�q�{X1������yf��Y�Jܙ@�O�I�PL=_b��7n�t���sh���<FC�/B���q���N�İa!oꁳԈ �RiVS�����-�k�{wS�����BAl<��v_ht��>�t�����8��VNmQ<mvMƜ��zOX-4c��Ku�w�+�N���}�::�wcI]G홭p���(��*n?ͨn����oz��E��?m�$ ol⠓c�~g�t�Ǵ�_#�{��w1�=x�@�M b=J����ɥ��Z9S�( m��?��ػ�oc���?T�y�r��,/�2?����D�e��G�)Z�8 �Ŋ�@�&h�Ĕ���|�tFR����W	���KȉC%O۱�������ǆ~�Ӂ��E�l�Useڇ�5�081N�kʮ'���'?�*��Qpb��_�fuub�Q#R%���9OVǩ�y�gHHIq���v"����$�4A^�)F�P{��B�?��K	wR��s}^�I�j������p|����v�1V�� �b��v��+�Y8�C��ROWޥ�y�[O$�5�5�k�Z$j�;�3���ʕ�2K>Q{Z�!��D�<�Q���4��%8�i0q^z�Es��r��R�d3�.���]�x���j~�i�B$��R��ᘈ���ʿ&��mi-�H# ͈"#��"=F3�F����Qҥ4�'ݍt�������zu�:?�7�#�����*�M���?T/����9�s�#v�Y�T�� ���A��vkr�,�2�W1O:��[���i�A�W!_��0f˒��R����{vcϽ���K$��)iy����j���(w\|I!�w��b�}7�'{Jv���$|W�ŉ4�rvPK0�y����������0H|�n[�֛���P=�N1�l�FX�7Ұ��vҍhl�ґ�T�� qg�B��%�_l�=�/���1u�ܖ5���2Сڃqf�VPa���O��-B����g��j���������7�$��m����C�W�}L�{������j�5�o.D9��N������I��l����[�9��Q��c�Y?`긟�i�{w���C����)�W�n�&�q����.p
.���;VM�VJ�bA"�*��%���[���쾲��vW���s����t�#�]�Ex9�ա]�	���r^��k�w<\��7���`���BE
���U�{>�n����/�*���D����?�����OvF�w��b�⣘|��ŧ@��(��GV�g��(Z�Ok]Gj
�1ՕZj��9<7���q������ �v��S����r"����#�Ι?e~�ڜ�"$����B�w�8HO_�W.�e�ў9X@��N����'�I&�4��B�Ǚ�O�]�X���6�h���+(�hm��ya��h�_�~���\0Km��u��ADp�y���/�_;���J4$qNr��2<�����h��)����H��B�'�.��;�brs��ζ@�N�2�z���`M�E�hL��d �(�p�d��E$�@z��"���������X�n��E�Ӟ��(R�Ց	�W�x�z���`Xȼ=�-��U.�� ����c���m�=	��Ǌ$�1�.p����ب1�"Iy��u�xo�������ҙÈ�1��tDB`w�T���a�u_Ư,��h��i~f�;�xǢ �l�r�L��Ƌ�3���T��V>=:��y����\��p��/�DnC��g�����y���r�����Ϯߑ��`N� ����p���kg�����M�v���΋�b��荎�'��R��~~ī4_E�)�~A����.�>�3R���l��t�o��/���g9���µ��H����t=�AE��~#�u�/`�:��v��D�\�C,NCW��~�֧*�ϒg�v]�}Db��茈���� 5�z_����;��|a������ۦG�1�1�m��/GJB�����`t�ح�[]������Ev��Ð��oMm �.�{k$�w�E@H�X��7_|��vۢ�IH7�{�E�ur��ڹ��N��iy�$7�	]����������Ӎ�!�����*���7;#�=22�tr�b��ތ���$>.t��Lj�:�"
n�ߞe�)��b��Ɨ��i�5��f��ڋ@�ʑ*s�}����~�z`��^$Ґ�G���s�TJ���-��7��iE�|�q�a�J��"Ph@k{��פ�G��]��9�g�TlL�UV6j�՝kr�Lы��C���T4�j�������!<�\�V�|ಗ�s{�;���LB�<���[�|x0����Z�Y�ص��yXz#d�(!��&�������)[�݉1~�wa�R4q��������s��G�H�_YjX˧wn`�9�Fʺ2�`Qa�v����U�������T�ofI�W�^1���	��N;��e=�u�
y���ͼ�Q����sx������xs�V����~�3�-6���v	�2��_,�'��S�Ȍ y�pw����ɠG�.W16��S��$6�W�:��FQF�>��Ynm�����*����n�F�b�~���������3��Dɗ�Q�ٚ.��+K���y�^΍���]佝X��$����dh}���4�=���%.��͙s�2�F��l���_
h�i�;�*p�<�˂�%�Ft�~aʇ�8�4E����hAQ�����9��G���}VS؜��E��8�v8�15�������	@�0����,4u���z��@7B?by��Nj<r���>��a� e�(xBB,�m���Y]�q��@�,#,�(�|�ÑSJ�]G�N	����t=�j6�S6�c ���fH�2�2FT�#Rهl�����b�W�
�����3�g
��GbW8�O��6>��?���ǧ�����r3�x�J�MHN^�����*&A��&���@�^�H�N@��`�6g�GhND_q����Et��9�\��[m��^�I�woח}�9ث'���� �u���cN�o�h�9����r�T� X�&j�5��~˟�7?/j�
�S[V��xL��J��,LD<o�@#�c8b��o�i!�_y§4f"�������Wx�'����"h~��gށ���ޙ�nH�`ycuE�� s�ٺQ�z����T�������C�"~U��,�'�_���>�{�d��r�1v���񏚩Utw���[�1��ߒx<!�ĥFZ��:�m�?��[�Cfu	ݫ�4V^hr�d�o{ұ])�W��wkf#��>H�ұ�9��J�fk���y�6F)c	����C��"�F�{����y�w�#6�$��>}��|�2&�����}�/�VÓ�#:��DK�|�.�	����װSӥq����՟ �`?�U<k�7�sҲ)t�6���	�_+��%��'0�F�d���q�J�_n6��,Sd.��k>�g�_s�_���r� �ל�lnY@�7E/���l��.:R��f�U�I�կ������Q_�9�hu��b-��A��n�\�l�Q����+�Ts��m��V~g�%����������%�#a�i./o������j�^+�D���'�{�f��$;dN�C��S�tL|�Ĥ;S\�N��)��W�g|��ޭk�&S-Q|SG�D�u�Z�9U&=�9�-(�fw��"��S���^V�?���_)!�'%�@/;x>o���x:>����"Q�F�q����ZC�Er��������R����J�a�7��V�?��N\�R0�1|�`�ئ�|��dv.��0��DS:�����5N;�B%��þ�c
��5�w����/�ӟ�c��3���E�繋V�8�2>��E�c��_
v�3��@҄�C6͎
9ڡ�o�7���:v
3S���a�z�(�Z����I��_R"1|5[WP�t���>��!p�ſ��H�Af������o%Kx�������������]:��h���ʂ���<������,]MΞ�C@�q	d]�-��T��Wɵ\#�!]����m$��1� S�	�ю?���
K��*�El��6��I���괇�q����đ����Y�D���_n$uŁO1���%����U�C�����uF�媬���E���jc�����^r��\_;S�Jh_�\j�7t��>�S0\{*�c�F��T���gl�9��N�rv���͒Es�_C�寤�X�����E����Q�_?+�ppd����P�!�6h��N���x�����$.�5'X�r>u4V��:�r��A�w �ȺǤ��gy=4�tʃ�	����91���m�9�&&�M�d�hp�CL�����T�ikcS�St�����m�X�C�L5qɨ��J�ʗ6�mv���ޗ,�<4)/hZ�ޠ@�I,�]�$ك���7@J��S~h���>���2{���d�na��}*����/[���0�J$k��:��&wgM$��LF����	�s��q
�!���e�I;k̭�H7��<g�1��)�O�W�����7M�J$�,��.�Jn_`�e��'M���B�J�;���p��;��Û�U�A���u⍹��퐙/-���_��}%��;~���8�����F���*�#'�æ_'�����D�^�a������TD���o��6 �I�NWB$�V����ƒ[ I�C��yc��.��_'3U��5�Uv4�m�g�m᥎Al�0D�~��hʠΟO�ѐ���n����/A��"9��r�#��.|C���阕,&-���⁐�%�s�J���B��&u�;��s���(��=�*�TU|ZA��@�ՐL�Փ������}�v��e�G�ؓ`�I�5��aw�3����liO��?ѷ3�M�Xӹ�!h}�1y��hx�~�e�x�X����.�	m� w�P��c���������Sy�S�:��Z��:���	��.���%@�!g\���09L|v��'~�2�ڨ/��<
S�m�*�M�D����h�`�_S�qs����8�3���m{ڸ\x"0��5��qϟT��o��|����=g�F��oH��<pq����&C7h�-��3�n����4Z�&g7�;��S�tÓ4)����B*�0bd�IvJ���,��̸���魑�w����!�~	/��1*4z[�\����I���.�����j��[]�W��]x�oZa�u���7�h�����I�~Nt-���ba�@�~��;J@c�g0�H
��B�����g>w���@�L蕟ч�=�Oo�^�#B���"�h�Y�)#fwRb��S_�Þ�b���G%�z�q��M�O�[�7:;�8 ���"8��<=k�q�>M덴���<��N��Y�M���l�߇HK�z������D�)+�PU�V-\yo����捯7��+�Wk���:>��	~�N&�V� QB���8��
��[[U��H%E��T�f�U��ME�
�x���O�(�J�y���7<�0<K�B�x}Q*�.�<��tۋ-i��q8d��pޝ�&��x�S�,��aZ����?�o�E�0�xoq}�A��D�:6uL����M���a�X�����ה��|z��]̛�P��!�o�"���v��X@b�xm?7Z��m�>�{EMQ�=�T���Ť5�j�C�&���$qoS!_4f[�����1���<���k0]�L�V^jʅpG>�r��,�%L�������1i�̟i�~���VSP�r�-y�؛՝.~a�/w��q�v�����0��1A�<7ope��?mY�?,~��I3�c"�lH����&�b���Y�_U�W�f�=I�Ҟ�O6,wH�:,��q\�;������c�3m��֛1�9�W�v4���X@���'�H,ZM�l��1���Ԩ=���{�z���.�}��pqS�oO��B�����vs��y'���Ys�i�7{�}$Rf�Db���j9�w���ܥ����I<)���s�A[�8vqR�3�\6�*^DR������/%e='R5#��W�}/v��%k2�Lmr���dc��k::�x���QU(�c{�Ʃ� ~�J2�?A6�,Ӂp,P���J��\��XH���۝�ru=�3zqq�UW�+����Y����g��.�j�I�$�O��U����+Zۀe���W ��O���]���lH�q���{�F�_��l��܏SoUPb)���N2w�����o�f���+���(Uad���Z�g��o�����i�]j����wOLC�������he_�!&ó�nҘ�{�Հ���gq��8$g����~����6h����Ԙ߇c\ u2+�%�ȸ��5颁�z�ݎ����������s��l��³+�pr�)򷸃��}Q��#{j8���~�����ɗ��LE\����"���C4H�YL�<twg{{ 5.ܖ�:�sm�`?J��^ѷF���	��V�iP@��|+�Bp��x�7$���Ι�v�W�+����
�<��9l]���x�h3I	ל_U�dx4of�ݕ��n/akÛY���H8�TcsC��O��������Uڣ�B���W9�F�#��.������ܶ�m
�mKF��jc�X-]Y���j���ҹ*� �{|7}m>s��,p�r��P	r�0x����Ҩt�:����|&-6�eR.wJW
�K^��v �XV���/�\9�R��Q�խ�J���U�+ye>#&e�S��&���	z��V�%��ڂ��6�D����"Eل4�����+#�CGZY����D��h,����Ё�����>U����.0eIz��:sjvV��
����rqQFW0�� h��; =��	wd�g}�>��='!6��-w�۬M�k�:"��R����jK(+-)�o�Ȳ��H}Oy,:���^*�YĖo��)�������M�nk�gp�Ѧ*�x�IJy�������n�%��������0�]��>h����w�wG���-}��ć~EC&׽�?���
�H�V~�Pp�KS~��3�N��찻�����y#���|8+��2�A3�
|��O��*��˂\?�T���J��;�ZZ�I�=�7�-�1\5)3v���fT˹A�'
>���V$#�$�{�<���l��-O�n A#C���
'4ȴLC�A�%y��V�+�|nm&`D�Y؊��b���P��E�ʬ)Nk���\V� ;-QA�\�Y�BL~"��`�/�L�-=tz2�{|�à-��9s��7�����p�<�;&�SU�]�h�e|9L���	�c*J�3�zqW��h��m9����P������Dͫ��Q`��A�Y=�b�].o�Q�Y��_�y�%kbK�_ˣ�ڰ҆�r}6�6��w��z �\<��PO}&Z�����\]v�5_�����ݼ�~[S�J9i���ʖ�C�2�M_�7��&||Cհ��u���k����Q�<a�T��Z�zU�$�
���G�h��h��Ǳƿ���nD��Q��;;/B*6t&\��9�z��:�uuT\�'2-�R4q�!i����k���w���}���)��`�%�K�X�Ѣz�X��6����ʂ�F�9ڋ����w"1򽾮���y���!6��{>�fY�g�n��#�ڮ�w�o��3�G��[^6����l*�ܱhJ�&��E�d���]m�G?0��(�δE:+<Zr�N�JEA"c���t��c��6M&L�oG�����$q�ȝ?��K��޳o��X��X�T����lK�����o'�T�t�r��ܚ����ʖ�D<�����<�ޜ�	��@�f��Gbx�]>�u4Δ��c��2�#(�1Wc�ߧt��VR`w�dգ$Go���&�%���IU�O��� �A�x�})o�W�a!B�Dl�����)Gcߔ��ň��S@�|i����m&�]��&s�A��R���Fb[RW�>�#��R_Z��Ju�9@F��j����|� �|��b��*.�ZE:������r5���8�<�Oٗ�QҪ�˸w3������QFM�H����d>HKF[)��2D9���6>ij ��r�+������e�x@������#bb/K4Q%��$����ŕ{��b~������p�ϐ�f�v-��;��mG^c�d�3ʚF���;�f�igv�&�-/>mb�\�q���-��[i�;ح`Vx'�_��ցE�⡡=��+J�0W���&���iqW�_���0�a��C�d�I����6�o��W�b�_��9�/�x�+�p�O2'�^)�ү�c}�d��3��n#�g�+Nne�L�qX~J�)�p���# �ߔ�X�M��)�V�ҩ;��M|�j�����/Λw����q�Z��-2ע�����$2#
�2EX��H~-� ��}�$g
I(Ȥ�-���	9��SZ�h����f�Zw�	V/��������#<1�j�?j��k�����LOS�+>�KF��b��ST�秤J/&W�=´DRNT�{���G\��p��8�%\�� �8�܎��1�QI��KpM�
l�6Ot�9��)����Ї�XЪ�~h������s;@dl����D��P��+qp�;�g��dA$�HͧuG_�1�ui�ȏ(���3f��\4���'�������]'���D|��r�u��s���]os#rd�<�]Z��eU���|O��4�,���[�y�R��r�����Tl����u���=f��V2�Fe_e�Jث��k�h�wBK͸��N�m���R�'A�hG��;9���*�r݊yF5��Ҽ�oȬ~��5��bV�B P������w��Ոл�cF/P=��(5�)��<��Jx��N�bXHq�j��$${���I���qڔ3���ic2�G�;]^�8�_I��[�eO���F�L��Uu�^QU���Q2մq�XT�L�-[j�����b=N9��/e�~�FI���(������l*����<�xg�g�Z̤t���9��3�w��ޠ�'�)����t@m�~(�?Ĭ�g������ư;�H���t��+���ty��v,�Щ2��<��g����sL�J��w.�`~-[p����UF�(����j{��y
�qX<�6�ǉ��?r� 8�H�� �s?
^J]����� �Ͱ��C!�Dƣ$SAV�c����M-<j�T���h��y{�8Tx��U��X�󌻿�O�,x�k0&��W���ώ�q6Z��^��Ή�����p�����6e�����z��H����������N.�Y{W�_rj{z�ΐu���Y�m�2���|��S�U��۝S��}��i`u[�������֯7�)Z~���S�I��?�P��c6K��W���޲ZR�f�r���2����"�2�}���,���K������Ɉ�E�ꔩm�b����׷)U�ܞz5�F2_����I�7Cʄ���`1�{c����l���Գ]��lR�E��iۥh����s�_��PO�ZF�.��\��O����Z���6�5�����\M�}MN�.�����H���u��.����F�_�;Swoy���_�c�ѿ34��5�TdKT���K� ��N���_�,������);���~�/�%������ ��������Ų��B�-�z���tks-����BE�R��PK   5^�X:u�� �� /   images/3d480ee1-e9cf-4ef6-9de8-5a7043d7f31b.pngL�UT]n������6���K��4��ڸ;AH����4`��>{_�1�j�����Q�t���1(0���UU�zpp�[pph(�WR�x>�/��z� ��Y�88:8U�����C��������ޯ���F�.���z|�TM�Xϔ[����$?u��@`%�7�Z.�c+<b,��x�I:�U~vB�������JAN~�3	y�f��l�g[�3���-	�'��䢻=��?/�fߊ��Ǵ�2�2^��/[��QG�jj���k���������Ȋ�r�ۅ���_���;�r�qY�d�>{4U��`��	w�eI +���|?�+��6�)AH�D����1l��]Q6��8���y�&R��zF'D�h̍��(;�a�/�����������}�6�'((�WX���GcM�����9έ#	P�I����"�=\�U��LRct���[��?���IE98L�)L���C�����#&��ȃ�qY���$��A@�K����'c#i����3��4S�Xa6�ECGAʯVP�#��H϶��n�`�,<}�5��ϖX��?���\�� eZ1\$f2�4Y�Fa���;�0g�y�X/��\�J���~m����.]"�<����1�)�k�l�Ѡ���_�-=@�!~�65�s�����q�.�Tڜz6�,-΃��L|\�4qE�$bV� ;�`p7���c�A�ƒ�N�-�����>>2���C8�>���2�O�h.��@��I�����NG�z�;*LVI�����(3ނ��me�����(�n���g�+���ռ��m��ni�n&+����N�5�;���~�.��$=��6�=��f�I�J�C��/S�}riD��S�	?C'��,>Z$@����Y���m�J�A2����-"�?�]1jZz���1lE[����{���=�8AX(�
���	;��^�|X}}�d������,��G�mf<7b�~y�;�Ɔw������8�4�Q���s�/M3-�O��\V�$���Po&0ۃ�D�� ��Ҁ�I�Onf(�_�Onw��0�s�� N�|�Ի�S���C���J���a�Η��`�OAP��ce{���䭞=�E��4�$���	l>�ehX[k9���@ݲ�X�',ȅ_���<�U���ٝ	����.�H �H�(���l^����+��`Ҍp�����-��G9Z���|�5	�܊UZ�C6�V�@|ُX��@3I�L��%��qes��^O�?0�K>��� �X�Ak��lh*h� 1v]��P,$~>��;ɮy/����h2l�y"�T��.���&�Cң�#/,
|[*��B����Ԁ� !
�ua�Tx� c2�y�
:�'�]�s��⏔��2:5���CVz�,|��ß�+���G
��~�����˅9븄��������v�A�H(ջL�
\�t���I��^�=4�}���x	��o�F�l��>�?���~�P�Ϗ��2�Nv�U#4Z�����<���5c���s�9t�m�{��X��b��.��]��0,����2
#E���,x��CI��MTHY�,��`{�������#���b����}ި��9��?�Pf>�I���
��������F�V�b��~��k�]���6��H�<O�g|�.�2���@A8&�ȉt9�kxRS9��_1��x���>�69K�{���K�����^:��3R푀I7�cD�<���Y�F�	�wk�����!��FY��� (��o9� 1�V�'��P��ڇ�>��p��O*n�ʞ�ik�a81��6*
(?�8�iV'5�<.��)Ha�hMRXxF��U�g|�7W��kt��"��J��_]�C�c�D�t�e?l� m>e<�_kT�3d	.���u��s"f*]��1��-�:ur��u
��4���A9��X��+��+�d�ڸ~,<S��xa䖃��IN���N"2��:��~�4����w� �������o�/T��V;�-�T<����xV��+�G�n應��D<[�|�[s&�H���"����r��A%�;����X�H���2g�
*.��N�YlY<r)�-;9>c���V���-3&q'`A��̉-�/��|��%��k�/$"�u�����}�j������e<��}O��q�kO��3�gVD��?V)p���i1ė����=�D�2�!�?
��U}A�D��:�g}������@�nz�|rT�"�B� ��X|Nj.ǂ���3lo�cQO�E�����BPP6=�&ⵔ�����?yT����N1��B4�^�Jo�������b1�%R���L���^��}����*kޖ6����a�?!լx�Ji		�4#t0�X_����������F�����L��R�n{�ۡ�����7�P1@��"^��6l�ŗ�#.��0u��8T�4�0K���u�I�?�#*$6��t��[���d��;��(�A�Ӗ:A�"i.E7���TVV��!G��5��y�q(�Uq�`�Y�l��6��\�%�L��eS
�'����m.���գ� |�e��\.�,�����?�(��K�Q�+]r��W*�?H��Ǭ;
P�A̡�	�Ob��&��x�	�'�b~U��`1Mj�=~<�kҕ�b>���ؗ����9�Ė�N�Ô2���>�����.'�K�
m��7�`(}h�j�f;�	o��HޓjPd6F��B�%(l�FS̔��8n�[Rc�d���p*�0t�"_"9I�����и��p�lZ�eǜ"-�+�*�p���
�3.D�#�x�/���Z�4�PNէ5�a.�q9����H��.�5\��:_�B���)��y��H7��Q�q�8$��L�e����ĶդSDr!��>$��ɁW��菢���`F��z�%S-P��XA�(�f36��� ]%�<V"�����K�dr����.H�L`�y~ńV�܌���b�C��j����c��agOo���d,���/�w�^Oh��	ko�z���)�8A&�N���ULR����:e,��7��F�M�[9���ƚ\�~�@�-���Ë��d=��s��(¨�F� Zga����e��0��Rs��ZA&�g��M���CcZ�:$��FR�(;":�G���N�n��˚���OH��Ks���;�2�E�X�Ĥ(�?58SdI ��/���t�
�(�'�]ܥ�pq���u�Z�G)�����"���w�4q�j�.�����!��i-܈�rcCi�T�g����L?-K&@}O�B������T�j���6%���QH*bdE��ɆC#h���a[���F
��҇$QS�P��a@���m�^«�ӬD��ԦM$�*��'���ŇP��A�xq*�h���T�R' ϐ�+5��#9=�N�1^6a�yv&���q���$ۢ@�:a�|�eH�D�%��3?���7��؂��G*�0KL��fL�B�р����?���F���G
4�=+%�Sp0#Ȝ!�!�7(T5ub���n:f�D�����@Y����ۜ���L��ot<q��A��� �G=�����Ac�8�r�ّ`=�ŗ!>d^n4|^��[�k�Yp����{�`վYj+GH!e_{y	�,�����%="��	y��T�%�i-	�f2���<�]�����#nSL܅�.m��X��7U��/�����a��b�TD`*��Y�{�b����H����7e�����2���,ar6�y��d�JC�a)gh�
yRw��+���d���P*�A(��P�
��T �8�!�*�	�-Ω���j��*��&$y�  y�!�@���D$�:�i� !����8t�E�T7N�d�MG�0%*���!�$���m�L�7[B���hl��1����6'�P��ĥ �f����65K$���&�H�t�PF��Ț�#t��n��8~<��A^0�r(����!�zzl6�^)�}F?h��r��D��o,.�)fɡ��Y7�^��6�i6�RUb���V--�(1�0��+�f�J�!��N��y�^([BZ����Fa��ɩ�t�<G t�*�yi,
/��b�aHǰ�n����U`�~4�CQoK��πo��g���V��`Ĥ6wFK�t�����h�����TS���[����X���J����M��z3�O�\cA4$�ػ.e�OZ
�����!�g9�oR�����pk�-.l7s4�W[z�Cw� a��h���)�RU��&�+FhL�6�b��G�D���/��H!E���O�qU����ٖ��t .:�v�g���L�j��x�c�db���5�?�����\����[EJ�xmل�I�8�"�p��T띈Z\�>�S��Y^�C��B~<޶]�0pc�)�R��WW�$�����R�V|d�R\����S�����ሺX�[[!�5��b�?�/�D�0���'W�)R:L	!��]@�H�tG+[5�
��q1�5.�����[]R�&(wB�
� Wn!W�a����Ĥ7|�5ΫI��l������A9D���l����q��/�"t��*�c1��B1��k{?��ڥ����H�_�����T���/�Y}Th/���ό���t�+'5�c�u�Kґ	�;��{�-�E��Jl�m����SE��y�a����؍����Y`ݠ�_S�J��`�!�9� {E98ܻ.�\^^��k��Ff�&���R���j���9^�G3�_k�@�B�H��ܿgt�������w
Eb���k��T�1���Dc聉�6m�;�t�2д�8�r�z�����d�H+�Ac��~`�6!�s��:��$V��|ԯ˟�����gw�$��S'|��~��:z�b
q�~4�H�	�ZyFne��6���t��>�3?����7��CW��xj��At�;��-��ů�l�T]*T��b��'�D�}8FZ�\)�e�M���p!o=���=^&|)�#N�U�LMRR��� f�!��j)�^Y��\EC�D)̎%����A�ė����ē��wC^��[�K����].�y?т�,񐬻�CGO,��z�/9e"�n{��$�y_��:1�A�D�U�8�{|EW��?O^ ��ď���M�K�e8h��͋��T_�l�Iks�~��*O����|xld��)�g��8�%�@��ֈ�icDU��F�{�Qri��sH�i�	,�+_e�Xe���r�KWԑ�A�#�`F��%X���D^D-겪��Om%v�?�X,�0u1�Jhy<�7����@�~חJ���
7��n��Dn����}��7��� ���͔DYV��O��1n�$9���5����bH|S�Tߘ?8!�-)�SJ�T�4a��Ǉ�?�hc2J��c���"�=�mO�0��b�J}P,"9��-=�х��ˏ`ч�1F��mPZ���
o)"��~Pc���KX�j�?�����mfsX�mqM�u�X��f�c��ʌ�N��(!�gԃ��T���1׮\��c�@JE~4�	�m"Y0�E$N�o	a��)���aw,K\�&���-�W_ٿ!*�@Y+��I��m%��⿧�5'����Ⴑr�
�~�x�a��l@<&m��AL"*�U@�j���֒쒙`5��:,��1���w�c�%�>��An-�S�#����IMjH?~ĺ��I�%��]��d��U���b�����,;}o���Bv�o��mR�����_��N�ΪK9Η�*y��"�2N;"C~B"�dN�qC��Cp���9��:�*1�1��� ��vuq'EF��~�/�@������=r~��;�����Q�4�� ��&CC��2�0��T�X�/R�f�I�����J/�&�Vͩ�Vv���t߹js0,tdG#�����mk�p��q�C��a^]�WK�|����"�n�JMRA���D����O�ĉ��܀���ET%�+I���@�6C�k��`�S`�Z�2jۆ��Ce��>�R�DA#]�?D�7{3�ͽ̤@Q������P���4]�YO=Z>*b������D�����k��X�P�sL�&i� h��X�͎�_Lb�"�Q�:�2��O��e�x	j&.��(�6�$W�/:x�xJ�_=<�#-E��O�&��ۙ2����k��O$��B����ǩ��M�z���Z�Y=z�� )���8�$�b7NY*�~V�UL�Q��O�ⶨR.� oUeuMG�O.j�[-b��qX<1�h�O|v�v4�·"+�e���{�I�*��S�s��֞��48��ȮL^�!�\�+ӄ~�-2q|� ל� %�\�M�Ŋ��Be�mce���d_3�ÕރD�M:3�!�4�iTR� �ӈڙ�jeD�QZ�<{�2pf��g�~�yȪuv�1��s��\?���si��=���>n� ��~��dE<&�*o�)�
�'.����7{��Y��y4=O�cٕ�=�C��.Ν�(�
�%-��i�Aсˎ��ʈ�kA�љ�»�wNß���=�@��1t����Fz�m�lQ�4�-�F�H��Z2�઱��*�T���c�$+M�l�>�h��H4�b�l.�x�tﶷ��}�:�"`���5��JP��4������6+��3�?�y��ىԠ���aF��(*�u��;=8�US>h(I�-}Ý�r�1P�0։�[�M�h�.�= �↼�V�Y ��y9,u ڡvZ�^Ȧ��d8\_d7{/G�.�'ד��`�à (�6�V�R��(����(�����ȶ�:�Nȡ�GBp��&7 �n�ꌢG��'��\PS%�WG0Ð>�QA 2�ԣ��C�#�#4g����#��$�v:{`t���,k�OD0O(u��Q�b�����j�FV��6���D\v���6N�7�<�A�a3�������QN�K:������H�����p�H��7U+���O���
	�^�����@xT�H-�����z^�
$��ԋ�S�9�,���K����F	��
�G] M���'��$c-���md��iP�4҃��y�/�����(X���Kd
�t���PS�ͽ���'�~����)��������:�C�dq�x�<�j����CY|�P��-�@�fu�u����C.6d[�w5������EN]� �F�&1��3�N����L͟&����B]�CXw0�����>07�x��7�Y�gL�Z��|󵝚��j=�nJ)ZU�@ٔ㷔~�Ď ����#���&��=x&�،��@g�r��'IQ��п���߅4Q��v�=؋�f��Cp,
�NF5g ����M������B<bt�=�W���0�f���2b�!��� ���������u��K�l�#����3&��5�-Z�����5���&;�bnV/�_��#�[�PS�U�Ym���	s�(�o � "H�)���������f%��� t��}yҐ���L����Gm�D�!9j#��Ԋ��ٻՖ6�Ĕ�6hB��`��S)�=ޢNk��do4�a��%�)Ę����������:���\�Ng������X	@��q�����
�t��}�zR�o��%�Ѫ>�ۍ��C�H�9nʐ���h��a-7s�<dKA�Y*��ֵk�p�p7P���x47����.����-�)���q��]�?pv�eV��ҕ�����%*����zN�l6dފ�?���e#gs$�y1�*��)�|C9�;�{�e'�i������S��:!�[Q����i�
�{�<�-�&a�[���͑�N.;�T3^g�n�l��jM��,v��֩N�n�t���׶�=�uoʌ�S�� %�^�8��d��CA�QX#Uru㢕��w3�T���p��r�0v##�F7�6y�&t".�If|�Uo�!�t���1��+Q�H����U��f��� nh#L�� ��x�z'��X��{�)�g����;�T\�y��c��Z�'��L=�Sŷ蜜�zD��;���1��7jE��UK�����V/�g[��!�����C�6��1���L�"u��k�'W��9 	YM+(���\i �͝�`Ū�` ��>��u���x�^��rP����.�e:�XL~��eF�G�0�0��Ѵ���F����Ʋd��`!%$M� cN	~Q6��4���I�!�~H�,�X�D�M�x
Һ���5�� $R|HG�@�+bӢ�)F��!�pfVz+�5��U�:�> F�uY��V�:E��0���Ro��{0W(��'�(f���*�x� h�=t:ǂ8�r"��2ژU_�8.إh�����!�w��zF�%C&�i�PK#�V��[�uY��O}��3�Ă��S��h�t���&+�`)��Du�_�){�����(��3uL<m���'J�Yy��x!����ō@{�S�e��)_�V��Q�p�Fn9B�x�PQ{���չ?�wasø����,Ԛ��G�N�ֺ�]��U�`zB��|����u�&���s���p��~�s�ң�ϛb�Դ����3%�ݭZAA"6����IM"j��K����j�e=�v('GÔ(��p�R�xG�NrP|�jI�pȯ#qoB@��ӶB�+�:�b�A<
/�~��q;�i�Λ8�~-K�82�tNԣ�#��FG�ӭ7��|o4��rO�h�}:#a��5��ih7e���fMu�r��l��X���F2����[d��<���%L���{Tl�F��M��9W����z�ſ~��r��4nK���
��nl�?��>,t��[����������ܫ�����2�|�'��sAآ�l�!�<A�,v� A�;$~an��ߎ/z�lNP��X-��lL)Hz��ПsN`/G�o��G!W��Vg,�.g#�줢�������]ȵ���8}t�{����#��l(�竮��wq�H|�5V����Qo����0e"V=�Lzf���]���P}��X��lܺ���LF9�ݡ��������V������
�D��f�%9��c
/��g�Oi�Ոﺜ׹I�b;z����-�<�d5�g\�ҶL�%L{1��Jq�
�P�OrF�NB#Ŏrhci֨�L����:��&W���W�0�c�h���*/�C1�R�&��U�%/E��>�K�%9�7
�xu�'�87 ��1�*�F��k�pԇ�C]�Ouy��0���7�oaO��N�J�r��"d��7h��
�gI%hDy��	P��`!^77������YH��
y�M-k���� �LW��4}�!��� b˗�m��^��sY�߿2��Cu��	�j�\�U�$�|�PA�k���R%�!�{/�D�tc�/[���SА��WQA+z#�t�qX�|��~�\7]���'�Gfe���xA�ZԚ�p'.�m�㇝Y2��J�#t4�5���W�6V���]"*��
�4�}u;�XR�yuf;��p9X�>i�������x��)K��EC]�ʍ�G��dXuO��5�W4�J/�4�z�ɢ�x���b9���7�<�R���1�\�]�N���&���!m�C��jyv��[� %}��&)g=?����I�>���&�#�Q���=��fF�!O��07��K�Z�8�h�YiS��#cq�/�4
���Z!w'�%����J���	yzfi�⸡а��Ȝ�5�D� ҇�>1j�2vaX���8.�L�,���EP��P���Ń��Q�n|���N�a5�G<A�G�D���N|3�b�皆��0�J��?�?�,�ZH%�b�\��� �~t*2��b��:Λ�zkoC"mo}L暹�o�>�7�tN��6`g7X��e�ח��9� Z&w�;m����ʄ$��z=pn��*�\����F��5��C
�̚��I�v�Ě�-���'yE�=������߼�f��������J�pQz�)�d���z�e*����P>�E?�Ky��֥�`��y)��58�Ӂ��dW#/�?��ܯw�a���Ia���+�A�#����=�ϙ�̮3����%&h/p�n�nw��'Q.���4H��J�BR�wF�7:C�D�l���#��	��/+�Y��r��(̴�#�4	�jD[g��9X�1�Py��B#*��;C�Xnmȟ%�7���I}uwMZYCJ���qCZ�JV�v��:�Tx�.���B�z��(�,t2C����F���7�\�J�]�l{Bś޽m19��EhBMG�U�T?V���y�����^2v���YQ�����`�D��[fV_�	��S�A������' e�˫8"/e]�y~N��o�L�8�k�!G>⤟\�>�8�XeYBG�zԚL�
�% 9����L0f�4�[s��[ӠI��U�s�D![E�O�F���co���s��tTX��}b�-�P��jv�ڤ�"�p"�+�#���aY4��w�(6~KN^rrHF�&a�j9�/Z��k�T6BT��j�Pt�����lR5��ޓZW!�=����O@j�K7��f}���"zD���/v�2� �+2}���8
Q)_l�fitd'Q�P"j��h��g\ʚn.���ڑ����U����8lcg��/��Ha�:dy*�Ϛ��boa���A�Z5 �;Y���?^�\{�*��ęvr�3%��Y��̧�w��yֺ�;��B�ލ���F��]�@���c�
M�j GѠ�7��̆��A��!u�b�-&�LWa[>����$�վ�0����ۥ�MիF�o�����έ�M�?c����;*D�]�>��n!�n��tlQ����7k�H|oWwu�%%�(h�C$y+�ܔ�%r΀�pe\�����ļU�r���0��@gm�.��J��b�m>� ��B�V�jѹ�eG[���M�IuSD=�b�\*�*�D�tWZ�cM�U�~�W�X���t�.t�����*y�@�sYt>2Ъ��@[��Gk8�_l7�����ˁnq��!��1�D�U q�u,�|�c�8�ZWFv��o�3����ȼ+%�7�LZ� }���.
��:�0�P=ym?4F���w�nc�eH-����A��1&���Vc��hE[^��x���t��ݜ��7�V�?3�7������KO��p�Ml����8�+ҥȿ�u��p{v�x'�b
�9�=Hl[1��	)m�;�c�I��F�]Px�g�?۫~�����	�0�������9`����`PB�α|n>��%$�`��D�:�b�_�GXe�{V�W8-*�T7S��isk�r�=�X�n�6+n�x���8�'������A�W%��Kߏ`���`}�G�|RtH�o�Ԑ��]�^G|a�3`٣ ����~;/}���;���R�H����� ��8@��.r]���g[�+��x��2R�-S��_�=��C�T
��F�����"�D12�8��ᕾ��:^MV�"�ce$S6�i��(J�};�e�^��bx�^���dgp3t����ޖHEHa�nC
�i��Ku��R��*$;�3ε��_M��t����bw�e��Q<wƃ�o!E�,?��î�?�$��|��f �S����Ǎa3o��x{��bc�&y�1�6�+Q�r:�DǽzZN�����;�L���Y�d)	�y�������bɟ��kuć 0�隺��<������G!��U*��὞�rF�� �f:���;�����i7$|4��Nɶ L��}�2��G#M�3��b������)�"'��EM��C�TW/�$��Hk�a�d�g58�2��>^����-�xz6�l �7����oq];�N�<ڻ�F��E�A(a�	��+�}�v�������ET*��C"'�h$F�7[�
/4;��4���Ѽ�jBb#6H�M*6�ޝ�hl(-�$���G<��@m�qGc�����3��s�x�8(/4Q�bG��#�>p��3E�ۊj�d�)�
p��-2�b�}gg��@�E�����!͎?"�4Z�Ua}qj��(�U��i%N^
tڈM����>ou���?YYKQ	���[�-X�m���\EH�@�ҽ�Ԩg���ҤI꤫銥1�6��zǥzt>��ªG�$�B�'�΍ϾKFҝC"�K���{	��J{���ѻv��H��|
�+г�К.׭�0d�LG#����y$C�(�%�ǖ,��^���Km��ۚ�Ŕ\����q��� �Z�M�TYFj��C�O_'����q� �sf$S)�;m� �sZ��ө�T�m�VO�^����Yșdu��r���t�����3H��(����h/P���ۚ�l�z
�lc��l�M���W��z8?��~5�u�a���)⫵�u5�C_��4��M,�:�F�j3@'8i�7�5����Ǆ��-z���.��V4E�gV?-���{8�m���C��2�A�Ճ/��T88�d�q8X)4 (��i�P��hQ5:�^v�/��c���52�{��f��.�c��_r��u�Y��j큉,�\"��C<�2S����)��WI�A�6kW�T�O�$aQ�+gT��j����v�	{�18 ���ҽE�M�FCD�s>}������i)�������:��)������A\gY*[s�����kO�?j�^~Ճ�:���V��6V	i<����>�	Oż1������@�Aӫn�O�)Z!�SZ�V����zO�f��T׺6ֵ'U������7_XK�1X�ǎߪ�I����9|�R�K��Q�a�1"���6�V�	��X�����7��}��<M��zS�Q`Mr����u	׵��� ,�+�_=�A�h�U$A�0D{~O��x�t��#�v�ջ����3�����ӇO0�mhB/�A�0�zG"�/L+������h3y`�ˢ����OD�k�
�]�r/hZ��rB����>u�:���J("���ELZz�C'A�-�^_f�
F��a�o-ڿ�OYG.�O�[�X[^̸��d"��ȩ�kWWlNRp�jI���E����19�,U���8@�8c�����>_�B�6L���s(�
Cѫ�\lmC(S�(����m�?����ʷi�l[鍐���}�1��,G����+'���%��3�E8��m�C�Q�zo:<�wpF>�-]��@�78���@�
�1F+;|��~0�Y��
7�����8�3e�H#�Z
��ǾS�D���{���
����vͬ���j��� �33F��βQ����s��/�s�9����¨��e#�mg4������*��VA�*�p�/D��`T��E��Eb�|%�C)�Eęv�r-�_e�V{��5�6o������'Ad�P��"oH�M�Y/��M��
u��O�7B���������o�A�Մ��z�n����;�a3Y�^]/�,��������.�D�C�����җ�� 
��4}X��$�{}��z��;fo��;��);kW�� �BQջ?uj�ZG0�s!2����j�L���	���z	�r
�������3�!�2�-�m��/�,҂ɡ<�v�N�t�"S5�K��T�@�a�K��n�C�!s�#���b�A�=N&;��&�?r)kRč��	��:^�so�������v�h���r�V��.F�~�������an2V#�'/�0�k��:����Ɗ5����)��ko����W���l��N(�]�N��Pf8�ɩ;�=_R�珠�5i��ȃL����w6��l_=�bw�=���6Z~���㖛D��*��fO131
)���S��à��}w�i=�=ӑ��K��xc���Kӳ&Y��t�P��{�� j�gVp�f5�����M1֠	�}�6�+�Un2��J���q4x.B���:���j�5D�\�aY<Q���!ט�(&J�)���s�%���:m����`4ͪݕD����9r6g�,84���D�
��������Pv�@�A~ݘ��2�Js0�����:���U�9Zm,Si\�I�g�����&�ђh�`����}N��JԂT#�����>���M3�|{&Ã{�t��cA�K9,"
j�y�i��a���l9~8��#�7�G�s�c�uo�u�k����{�ϘO7
SIX[W�������I�X]<�g!2�0�4��*P�Y� r�ʽ�r/�g_��O<���d_ڈ7�~�`ϋ���u��§G��;���)������{�~��dj�]�m���i�pzgC}W�4������Ŷ�+��M��4@�X�b�BU��R�9����[l<�[���{�j���1A���8|^
1=O�n���Н�7��G���� �$�{��_�j�3�t
�H��kq�[�ԉ���r@�'$�t�F�d�����\�v�O�>�q���C ՅE$�,�A��~	,
/e����7[��Q�>�C� �;1'�&�[51+��F����3iؕS�z)*�5���q���Dv5F�0�\�q:N�Y�/�uV##���e��{��_=�;�l,���"�;B��i+�J#d~{���5�5��@��i�3	�9��ԅ�=$/
߫ �K8-X8n�%e��n}���*t��"0�14���L����l{������-�G����TK$�jO��.�G̪7eX¿ix|�	A�*���F[*�P��o�F���hm�a�k�3�������gAQx~?}�x9z�_���2�O˲��h*��)7?A7i��V���ٍ0@�T��k�\��&�:�"�]�'�b�[[�9.�M�u����]�e�=��pO bߞ
�rW��;�D�\Ҁ:&��P;���N���S�J�
�:ٺ�΍lܧgN,�Pfci��"He�DR.�J���[�DcS_;�)䵀=V��&���/TD���2E����?I���t$LU����{���P�jonj�	����J����%y�
���K����H:p���\9<�[�#�'��)3���оЋ�c��3��nj��%���{kI��B�M�;�v��υ�\���88e�G�F
�x�H�����g��z�q���]�����&�ew�β�D��!��-_׿�����G	��4UE�5�Hy-�
��'��̄����B~iNY������'����u��U2���mJy���N|��ҭܐ�Q��Y�tY����ÊQ��ac�6�0UY�M5��;�4H��N��u�e�|o��J9�(��`Kh��[4g����Q���
��S>�O(����C�=ʸ#G�T�A��&�.�{��WxtH6i�'�^�r��^�t��e�9H��F�e|آ:C\gp�	-�A?^⺷�n�D?Jٴ�#�_8��?�5o;~���-�'���*�_OY����?�6:B��U�U���P�8T�(�022�Il�ٷ�j�j��������x�@~)!4�Й��������^P�p�Z\}��ɝ�8/}Q�n���_oQ$'i�}Z����E˱����)�\R�G�p�ԣ3|t�߇9|�s���38���ٔ�Ra�aW���)`�l��nӃ)�{��E�������D(��(a��lLa��!F�G�?���F�KXaz���9Mg:v�|�o� �V,�����-�^]a���[.��wc��eؿ���A�ǖm�Ă9R8"����y�B:��\�S=�&cc�8�NT�y��S,F���xD�����8A��Y���ّ?�	�'<ﺀ�a���4�;��FE~�8�F��j���wmM�+����#��a����Q�����z����)�fxTs���YA_a�h�i_9A�v!^��N�!
��(�Q����^}.��W�h�sT��w�α5�Xi1r��LE�gŦ��k��a��^a�U�lя�Q������4N��6h�/�8@��/N��ч�q���~��8�"%ovz�=�Eu�O��|�vn��:mJ
�9
�\Y��n\����=*����h� ?V��Ir[x�7��@]����sC''���֔��wgNA'���m:7��ȷz�o?\�	��e�'��,��pM�8�i8։_�k�;9�ɻ��P�0����P�7��>�ɵ� K���`^����^1���g���k����/�$5��H�kq��ji�:�kȭ�������<�����w��Wt��9կ~W��W]d�b�s�Pg݃�uqp"Ny����^�@S9��U�&�,��O<��o��&([x,f��^�ح�R9��R@����<#��5�D�y�g��z�"D�v�J�\��@���yZGN��)x��	F�!��x�N�esw�"3��/m A�Ҙ��f�T"Hp�/� �I� �Q��8S�fqq�o�J��%N���K��xj?��?�/�v��CM�1[��,�X{���!
Z	5��v�aF�a�c|x����M
.�X���	�Zn��ʝ��",� ����!�6�w�4���@z�o���6H�qk�a���A/�:t�\��1b����&._�����.�_l�ݬs#��޹	9/�T/aay�k<i;>�t tcR�ܹx�u3�d��<���G�dʛ��S<��(����&���e�w��9�~�Ӆa�0w6Q3r(�氹��8�A.h��+0����Db���2�I������v?���8�X�F�-\��7p��7����4�Fm!3�{�T�I�3�67v����=x��
�a=��ZF�/ϡ��>/}&ޏWN_�Ƌ�xi��3�r�龰?��7:`NF���)�;oZnr$BLRR�%0PS�	�yL ��Il�NB;��i���6�WA���fA�r"�mt�e\��q��_�����+mkǡf�t��s����x��Ӵ�a"|����/EJV?
�|_V���T
G�zh���@
OWȠ�Ê�V0)ħ�㩹*S�_ ��#�����)�W�^@7�^�f��o`f���W 
�5`��H�K[y��T��MCʹOp��3H�R�*:����ҥU�n"��^�S�K.
�x�os��Cॺp��I���%�|�M*w�8J��������%N���K��xj�;���N�[y���BÓ}t��Y�(@�L��E��<9���L���S ���[W )���eD�Yn~��u�cx�=$��!�a�v:v�W�_�/~��p�W�i�m�/�ܜQ��SH�"��*�g�Y �j(l[��x�������4�UL,��6dCbטop�}�R����P��s�H���z�5D?���v�R��'��2�<�5��g���	�	��*���G�7�*P���
����
��zk��X�Ǫ�"��2�媷ZH�58�̥-���z���軐�	�N�Ϟ۰�����m\Z�Y�+��K=~\�9��O6����#�C�%&1*��-��\_E�Z�ń�*l�"0a:�ѤF�goV�MU1��yśA�fX�O��!HnQ/���/;�-���א�\��#?n䦊�^;�R5R���N�ť*���I�}�s�C�c�F��^����;�&��.j���]	�9G�����}�����,�LZj1����{���3=�9�r��ᆾ�7M`�@.�p���(�e+�!�a��Æ �0���-��a6,�a�VZI^H�ĴKr�!'s�ܹ�o�PՕO�s��}���t�rwd� $g���
�N�����y�waN�U��xGl�1�f������2>,�֦�-�*K����JfГ����#���FcfJ��Z���Wj�T��A����ݜt!����^�Ǆ�`���- �Z��Aο/b�q�?�>���`i�
\� mf��:����Q/�.+%*��� /�)I`�a!��ҥ53���C�vɵ/���x~oo_���T]���M��A*�E�2�e����b̜���x�����o����b}����m��xE������(;��F9���*���A��X��w*�ɕq��@���������>FH�^�
7a�Qc�i��VP}�	`��p�� |	������c�x�?�\�g��j���GJ��f�m:1�mJ��֘�\Fg2Ҍ�]��͛��j���_���!�gfq|r<ޥ�K�?7/7g���5^��+eS��ࢆb�B2�����!���~�e�\�����`ay�Gm�"
1���De�W��}�έ���.�N��T	Œ�:ӹ�8��ڜ����^��w�:�� �I?��7�����_����e�����f�$	ݾ��;o��+Ͻ(/��h>Y�_����.]_Gm�.��򔦬���x��<==�b�0�X�'v��8�*5�z��S)@�V�.�!�QqNpoD���	Ey^���kG��w1�)�f?}��w�����̠?��s���D���
T\fPz
xun'��+�vZ�q�K�uG)��g��*�x9�ɲ�-�Z ����b[��-=ֳ��WF���"Y�aL5��펁�DB���f�^��_���Q*�%����H軃$xͣ� �ߖo?�`�5���V/�<���w+����O�U���S��d�k/9u�	�{�R���ǥe���R�B*�K��{{��e�J�I2��h�z�|��k� M��W_}�?��������9��~�f4�&�f�Gf��x�����͛7�����ֹ��L���Qvp�s_!�ݼ[Ǵ_�F���P�wp����(�ۘµ�]���1��,0w�Ge����%D��Qr�`�{�E�u?�\�I<�����9��F��)��p�Mq�T�(�h7;(��f�P`�Eؼ}[t}����0�xw���ħ�Wt�zi+3�U��5���p�Ow0��ٕ��2M�و��DY�o��;o��b�A�wg0���V�9�{��\�Ts�q1;��M�d�B��\>�[ȡ����������������'߆㟠�x�F��1\��%��3��cQ��g�� �LעL�A����m�{��D�a'����z�ޝ[���\��]D}fJ� d#^���ycd����+cW�����=����p�l��v"�T�E#!�	I&��q��Ocj2��p��-4���}˃�5R�������[@�&����x��G)޽_�0�������>�e^���/��;}a5�<!�ײ��N���xE6�D�����خ�|�����l�]��5���M5x��c^��:KY�e�)�3�%We4HR��\,$+��4&=*��	�
wQ�8hE�۟F��� ���U伪 /�x�JsH�x����>Iu<��S{}��t�T��'��wd��8G��V2�E��Z̝��,��:9A��{��=�f1�g����>*}�/��"�|��:���:E����76���3Ez1��r��8�
�B1��rS�^��n�s�N����I�Z=�����=t��4�?��x?�Kx󭷮������h�):��>�&rn�=���/V���bw��.����t��33���5�u��3=�t~�k� ���MD��c���I��n��cps����6�J�D�y0�\d0����~I��b���IOӾ	�C�8�M���9���Źyܾ}��ܧ�\�[_��2��@�H1��$$�tY�e����%�j���^
��\��x��(�FC1��sKh�t�"/�����P�1ؼ�b�bv�<6��э�K H1=]�_(���wf�\	q�G�b�.�F��Y���q����;z�Y�w�qq�$Iz�uxuj�0S�	�j�wwG���ﾄ� B����an����iT�˸x�����5mIi:^4F4�
���K#k{(��22�o���)��!�/�4�Q�u����Kcxi��L0���+�'�C�d����� 8��2����e�7�����ܯ r���_���9��E�$u���/��	�;��S��}�l'�r�Pd~�Рtb6�L�L�+���x�/���v��'��m0��v�j���QR���@x�>4���1~���'��������>J��(Tt�e�ݫ)�=����㈗�fF��..��2�=��.x��:=$�E/���9u��T"^f��e��8�.(�b��u��X)N/�#\/�Yt>?���~���ǓO<���F��S�ykk��_����w�OZ%?�g����'Ly�b���^Q����gggmm�? S�c�ُ���,/�[���׿��?���($}$AK����)8i��<��f���ҽ����:h����x�*����rf��J������U��?�(���0­]��I��(���ob�v�3r)����݃F�r�� /A�Mc��ߙĸ�6��.^���(��X\\�b����"ɥ�p�f��+[ʗN/#[
��d�' �B��^y�PT�{���r z�����SH��1��^��^\�R�{�(������#�-^����Q�n�Ӎ�Lܩ,���=� _`)�8x�M�x�G�F��ˈD��/�"�ן���u�X�ų^-���I;N� vq��&�}�~�e8����,L�Vs�����*�g�%
��蘾P��3�U�x��	)�!�Ͳ��L`=>�G<
�<R�Y�|a_�,�� /��ޞ|�����ߑ��L(r$%l�7y.^�px^����7��H����_��}� ��(q3�+����x��f�?'��X[�����!�R2r��T��1�\���^!�^�����Wg�
h�Ia��}����3$Wx��Q��u�ެd�6`i<��0�cDH�J�z!��t�&��uT����j�k�>�C�|+����5�xPxy�x�I�Y�c�C$���@�Gl�3/�����Ø%�����2;��ǈ��4F���W�&�vssSX�L�3���?.���/���S��?�t:�����淣Q|�C@a ����?��B�$�GzX���0�c��7H������8R��P<>��2s����?�Ͽ�7>��uTr1�~Ѱ���,J���p1fٳ�y�;���6�A�d���U�_��č0���斐6��]�
���&��U��� �F{0�{��iD�Cx��D�~QjA2�� o�{�F���N�;�U*���*�¥#�޻���#����P/ձ����_}O?�4F~���3W����BY��)fޘg����Ű�V#�x	����K#z��Pȹ�=I���/��(}�g�n���dw~cz~��{r�H��p���8竈>�� A�����?�x�O��ڗ�^�g�ɳ%&��Se���	���LO������D���9̽1?�b-�\���l'�[��9G���s�T3Y�x�e��L�1�6���@1�#N���pO�I��#6U�
�\�܆I`+L0D���}W�d��N�X�T��!��o�w_� �?�b�0ƽ�)8��0����r���K�=?�HF�\���$�#���u�u���s �o��\+��c*�*G�����U�g=� ��x����[�ig!��C�A�*F�+i��?��"^�!�>^��ϔ��:2� Q�G�t���*\�N���;��@���������X����р#^ac��ד�"M5��b�7���J�X����\G1{�����5�,hN���
rt�N�*�A^ׅ�0���P�w{{[�f���=Nv�K/�$
u�\���?��G��_�Շ��o��Ɉ�� 3a�f��h�{�N�*��}�m...~�����پ� �o�z���������x��'�,��GN$���Π\�����fS�­����ܽ��A}'���.\� �i��3�L�S�ȓ�x��uăo �n�������SG����~��9ʾ*�:�[PĽ��V#�����'���@��ԏ�������V�������3��/_@m��wxY��EjS�6�e{�eHJtg��R*���#ℽ;���[���s]L�0ռ�>�c�Y����*�p^�>���;l�q#x0K�KI5�f�#*T1�+�j�y��z��^}��.�Uk_ƥu���7���OL�m�#lo�`���z�M��|ו��1[G���s�sR{&��b�k�s�A_'��`25���Ff�`��K#��xً;�����(�+%�J�/(��(�Ij��
I�Ӵth&KQ�,W�K��b	����p��`_�\�=�o#���-��9��u؀W~3�?���Ϡ��T�0f���aJK[�B��$�zC^���}9�j�,o��/��6n#^��-�e|��#lm��a��k<~�,�����ӟ�>K(��(�g�UY�M��� n7bu�Z�?z��-8[��Q�y��9l���1��9�άI��#m�������B[�<�:F�(���"�����/J�c���L��g*�X	�\,�9Q�S͡ .��稆fE^������@L_{�����˿$�dʌr���2����xQm�¹s�L��p�֍`uu�KW�\��`�,7��~ �������W���?�m{��/��0�Q/�P����*XZ�����y�dw��1�[�q�1p���:�/����(�8�X� �"�=J�B~��{8�6qss���4�������TmY��<ߌcc�4���G�M�G�*k�	�����b��6v�n������"ί�Ƿ��,~��� t"�]���tn��%���˔!�����x>*���iM8��)�D�L�	�]����(�RA_<뙹y���V<��T��摤�k�E��n�OVoF�
ĞT��1��Q���{JC�o ���f�Y8ޱ��e���.}�.}3�K�f�uLrkw�+�朙R��<㐼�`w� ��;x��wP�
4�<�f�2֎�|f��j&sY� RM����^���/�UZBF�1�(�$H�]�婢BD��Z)��/��Ȣf^,j$̱���6pW�O��wQ�0�Tsx���m��68�~�0���Y�ʟ��◰v�Ө��jU$ӯ�Ӱ�)`&`�Fr�Q�h5�9��ݝ��̖�|�������U�V��'���̨�#�VFV��m�6[�/���ڝ�x��b>���˭j�����@ۮ4NA;�`���C�A����ֻ(�!�M
{(O�x��<��_�f��<}�[��6� �8�疤��t3�k�L�3�%����/!TG$Hr�FN�=�V��U�k�(�=�q��N��\>/ j#^΂&��K���5\R���"�A��k�/�����]�cR+>��P�����(���z1����d{�BIx%�~Gdi/^���~��?� ���&?�\�{��t�p&�����B�Z__o�_�������~���������RC���5�x��V��2���`�y��m��#�7���ll��#W?D���;u�3��4�d��z��>���zo�hx��ou�/}��e<��[���������u�Vg��[�b�� 3�Ut;�7��s���ml����^���������)~��h����1�4#7k��1��ޖT�;��sRߡ!,���=�����]�\e�25 R����7�z$�M�ј����5[���yn���قh��I�uw_k�E�銨W���pH<g�z�o�+�E�*��)�x��6��\��ױ��Y�/\�a�2L<�Ɉ�>�T��>U
�G�Gy��]���<JŢ�|	���]��}��k��9��c9�����KXϾ>�z�jzxmK�(Tɼ`v�P�����CģHX��2Ph��kB�g7u�DGG��������|�MU�(0�N���ڨ��'�1rv��[p��*=B�l��k��Py3��������*����8&��� t��?G�ͱ%��ڭ6�>�aMǡV-��C*�²��%��$�v�C!\���Z����H��u<n�a�}�4����{qw���HKOe)%�Ϲ�.�U��9������K��x�4��pk^� hc�?�q�\��C��>
^n��Y�'1��)T90��#����� ����g��fڗ��s\�!�8�t3,O�[�%��kqh�����>��6
�2�gg䞵�$�,3X"g���3�C�+�-9T�y�V�#����u\�z� �X$��T8������B:X�>�����/����������K�� v�#�͜ԃ��������7���;��L�a���4S������K��{�\(�]o�_���/F��e��Qc��$���f��+�o��§7��q��m��    IDAT�=黛Y��r���5��.�v���(���h�'}�eT�^�꣗�p�l��4_�W�Q��\���M�Ns��8h��ft���(��0����OE�߅w7�ߨ`������a��=A�^F��c�㿜6o��νm���X^X�ׯ|�+x��������ņ܌�"�簵���` l~qAnP	�!or�/0����C4�5 $㸋�woyd���83?'�f�nu?���J)hw���V>8�����rϗ}L�TP�P����E���$i��.�r�;�7�x=�i��wI0��+�~˟���e�3�XA����,�d���'L��8@�n�n{;��H[��55N"@0m.Qx�'��*�4�����-�x��R�Z&�oA7Ǚ��!v���g�x����}�KL���L�Jz��KGIF�%����%	ԩl�Q��������=A��#`땎��v��(WS��8h_@��8ӏ���ǑzU��r0-!*I�b�I!��4pr�
�CD��`(�O�6�&��=3��K��/L]�}��8�i*ue��=;��z�zS�w�3-E�1U����2f#儂�%���2T^�~X���?��/��]��' � �!�j����G��
¤�N1_�N����ի�M7��2N�2�"�9�E�*�E� �"
9��d�Q4�gk�d���FꕊN�b���͵ȵck�:���ZU"Y[��9�9	��9�S՚���9q=Y�\�G'G"��#ԧ�z��;��B�����$��u��~I��\�y�C�h��&�*�o}������q?���x�e���\}��W�8qݏ�0�-���޻7�u�D�T#�0U�/,tWWVzΝo-/�������z�\oЙ������n��*���b� 8�6�~WH.Ӌ+��f�4w�q�V��B�x=o{�������×�H��/#-Wx/D��.�V�gt�{/����5Oc\�g?�7�/4x�թ�IV'�!�V������(1]�3�pw�o��+/����4y�Q|�Ͼ�O>�	�dV�/aa��U�%�w��}t{=I͒��z��W3uT��MKq��Դ4���<�)�T�sIagLux	Z��`��u�r�{����Q�E��bz����1�D��P�P���PvP� D���I����� �o�8u nEN�����.m�2V?�z㲈���p�3bo���s�<h�٧Is�2e��<>��4��F�DEY��p�x)g)ѓ��&�q:*l)�"�^�7�>�Ѱ�sI�����K��ib�(r��;�X�rEU�M����}���BNK�.\/B<�y��`N���T^q��B������}��B哨U���Ǒ����d���ȕ�n��>q��� S<$�eE�F�#9fz�]��]��GN��:t<�����ű��c��'�O���D�g4K��66^ِl��0���8X� N�Cs�ԍG"cI�E�!Y�ܶ�r�"�2H^r#�N�4�sy�?��Ǝ�c��C ���Y��`�0���:"o��֦0�F�D�H������r�TjzOyJX�O�!1,��d�� �AT;�J���J}��O�g���42���Le��$���(�g0�|sS�Uz��7k�A��W�L7���9���	ח���A�q�l�uZ��&�&?��t:���b?��_��g>�aa6�Ƣ������֍w~��C��'���SʣQO6'���Y��a���O�.��Yȣ�k�_�C�|�e<zy�~
?�"t1��L/�X�cya���'x��ȵ��k�;�h����ױ|}n�NՂ\�l}w��`+�$c������Z�<�Q�?� ����U�^M�{���c>��C�~�A�� #Ô[��r���$<��믾�j�"-�z�[ظ�9��95hIIB�bE��oo�ddɴ/a�"M����V��P(<*����ޮD:a��`�L� 8i�ľнC�1�aS���Ĩ�+��
>���~���8<>D���;A��B�q�p(��u�{'Do`��3X9��(O�����U0a�r�
�t`�F�D{e-�Ұ�� N	����^dc��)?�.��e���N݊�4�X���������3'q�2*f��K c����/)E��yd֫5JK�Z{��J*��	�N$z���n��-T}��X���9�!���T���O�/6 ?��ij2nCIȪw	E���Ԍ\�wC�I7#QP�# ��{hLϠ?�HR�U~E�{�l�<��7�GP<D�̑�2�*ck���~WD61r-�3��|�I#�ֵ��@�sDp�}�����(���yf2O��r$��n,�)��aș�Lӟ��(�:�J=�JjW��yƇ�Ea8��ΣR�BDau7�0J��N�fW��T�5�����K���C<�c�iZY��SU�|l�{����'S��%�@$;�$���$ŋé[�D��n����n*pK������p�e��+h�O�:aWA���g�Q�ő� ��N�e+��I���r�>�Ao����/}�s���̜�X���;��j��������$��SO���q�#v KZ�|�ۗ�t4�x���u�.��O� wn� _x�Q��6
� �P��
�)xN+��p�C����(��"�w�H���v��.�zԓM��I��A��я��vu�nas����A���/!�/�ᇿ�eXgv�T���#ؒ�RE��oF�$HQ)P 8>hbks��4�S������s�`���Jv�Dd��
l�l됄(��@��x�W�fs�#�>��H ����L���tt�o��	�H��������
A�����5Fu��hً�av�� �s���C�s� -T�"Tg�pˇ@)F�-��v�8�,Sb�־�ru���l�X���&=�qz�6RR~*�(Q}�lYF�2��ω�_"AN"��D\<�X�&Sz<V:65����3mM�����x��#�e�$k|�haM�#�ث#f�&�U��#��g:�I����y�!8윬�4�2U8
p�i�� r[���b#�~~�~R��;N�Y8�*.�=�JmN./�lciv!娈R�*�f1��<���=8I���&�Dk���:5��(>�e���4[�f��-���� �f[~�^�����y'۶��`��vv�p��Hm��S����:9F����Wk���'Az��0u;���@�,\�N�����I���������R9/�`i�A^��L���X�P�JP(�(UjHӒd��""�-X98>S��A��06:����$le:�<�t�R�u����k�JBc%��-u�m��֯���\m3����2�\���a6�틠F��A0Q�U��'�>aϗ��g>�Y$)k�O���@B����%���fZ��(�sx���j?��<~aq��_1��Xn�#�U���?����.������?/c����EK :�H�ɨ��a3&����x�-���ve���o|��y�<��%ԓ
	k>t;=8^	�s8���?B����p~�C�q��t�+��zuN�A��@!:���)$e*�qa��a��o"Ώ��������%ll|�<=���>֧|����^o�r�G4���9"��u��&�{���z�����f�rT.`aiA�������]���:$��yM��9�M�t�	4|O�`��'�a����}| �fkwt h['�T��;�; <:A	��K��lw��h�]�̑Y;��0�U�=F;:�ܪ��E��t�G�9��G�+(���/��XG�fK''�D�?@ЏEĞ�U�TA.�a�)���.�������J��ȉ�mӠL��-p�=	<T�Rg��5�˵2�����AMV*����']��#��XaJؗH�S�"1�<5� �:qF�J�YӬt$+�Z��=��P���D���N���D��?Dc� �8��"�9�؎p�-"jX\��be�bIf�r?nݼ�h�,@�[��J�+E@�}�'�e}H���x4�O�ϖ�(WU�Xf��E��c;=*W%�V9���J%[<���qS��7_�}*x�$/F�d�K]�' 1�����kZ%��k���|G���}֘KEDi$�ϒ�a�SIA�W�ȇIp�<3�M9�P.`���5�2	�#����2&�[���nQ$��ŵ�{�3�q͎�����fFd��x���?�dK�9 YY?+����� A��f;U�J:`��?�k	�t��(�eAHu�/�I�6GLj�Du��� ʬn��%�4��}�֧�-�����Sk��}(Z�>^�ݻ��W���������4��[f����7ޓ��� �|(�(�$Ȼn���^�:S�1^x���{8?_A5�Ï�"C���� X���b�b:�0<؁�����i��)̬o`��81�u�x��p �Q�W�y],^�������ƝcL7>�N��{��\���O�P�0��e$��`���{!>�L�1`�#��E���dr����x������ۨ�a���~I�d2u)?�:9���$N١qdڎ7,of�����0wUp%���`N:B��C���Pp<�lͽ=�$o�Pb�E��|�Qg=�G�m)�P�/���B� NC4�M4'hM,�50���F�Q����!���,�V�@���T��p�l��u�5���z�1�`{�4�6�]Q�a�+�ٴ�8,���9X2�o7�������.��X�p	�����r=p�3��F�C�/;�Ϲ�/-'�D��N�.!�r_"�.��H��Zo��C���5�Z&��#G�u}�`�$���z}�yFP�����)Q�>�q	pr����AI�`��L�C��	����D���5r:,��k#4��h�6�#�V1k��1�,#�HX�-I�R���t��s���u呶W赵J'�ڴ�����%�O&��>��R�c��r�����1�ڗ�*#���z��\�H���8v�C��fF��"9R�ˑ��Ȣmک^�줯�o�S*�!-E"6���$�ڶ,��H�
�ک�*��6�wÄe+O��	���)ݞ��^(�?�z� A�vB� �YݝΉD��t;X���׾�|ᩧ���+���2D�+ީ���{��=���<������'153�����!IP6���Y�9.��(i��p�wp~~	S���<���WZ��'������P���."&�w\���0
z���AZ�a��:.]�����{�P(�9�¯W�O���^.�d��@�so���J�!籼�0j�y�.+8>�`��H�M�D?�|,��
��=��J��Y��N�����8w�޻qK絲vX,�GC����5��ӑD�DǜkZ,��I��ݻw��k�����5�Sq�o�H�/"�_�҉щ��(���6�N�N��
��"�5ʒ�lu%:`���� `���8t��n8D;n���f�kpK#��A���$�I�����j�r���0��aͣ6��W�P���8�y�0dj�7��<.��x"HoH��v���l+*�j��V�����5^�n	VLAK�b�MC�ԈQ4c�L��{.��EN�"x�dn+��,Ј���@#fv��+����z!��� �^�G���n_���i�
�}*C�[�`0�4��F�Mi�	
L��c �۴�ީ��/��K-��b���En�s�m;��O���T+Y[l�"������v!�����-ۙ�bF��T+�e�Ӷ���O P�����rq�)��0eKRW"�_��ٹL���G�gM�}��jŬV���i�Q�ZɘQc��J� 8�+��g�!�IO�\W�����V*>�,���g�����aMV~���a8�k�5�P8�(k�6�5]>8���@�)�k��R���(��}��E��gK���D����_�g?�ߺta�w��1��rs/�͝�O�k����%<��Ϣ/}f�0����s�Dl��MC%���{���.-��Q���p�Bn4D���`�Q "D��)c*WG=_���st�^�D�F�4�eL-/����lwo�'7S/"7]����*��M�e���wol#_��������f%�Y�M����Ξ�	�F��Y��P%)�>UA��ł����B� #�b�����Ćx�ݛo�)S���Ψi,ތ���dŔ�:I7	�R#]���TCCD#@�$<$4���FR��(��Ȗ��U����d�b���#S'D�N6�\
��)g��8V�6��%�.+�FN��r-h�9x@��w�ɔ$�σD
�zb�u������&ƈQ�i��[N�A�Yf�.�k�K��G4�4"_���8B��kjy\�#�]R���j�N���e� ���Z̢9M3�2M�&�̆YO�+Y�iݖ���1�H�|bE`MZOE[�J�)a��5FG�H@�,+����������x:%S)��~�� 9W�<$�ѧL��e�s�Ly��������s�kŴ�c֏�����4׀y���Թ�3�2J$�s���ml���n�`D.�m��9���PF���&k��u3�38��.봒�����>�����)qb�p�Z[f-X�GN��2�$��ͣ��q��*��,�%�|)���f�: �w��mK�n7���.\�X[ ��j�ncfj����]��_]�|�C1��#�p���_��?�ʿ�]Z��x)gG��?�H�F��{^�L�A����z�V�a�RC��ī���a���tI�/Q/�i�p�^n���V�)'�#�g��r!R�F�@aQ�g�W��>�J#?� �!m��rS5)x��nρ_�F/o�j�&��ސ��(�XV�W�cgDT,�0tP+0�uA�G��F���L�B)޲Q]"�Q����.}�њ�!���Wք%�r���a�jk��k�F�Fxd����S�����2}�T�Z,�A�!E(Z�Xz�y^xň?$`W�[>�)��GL�H-`!P�Hz�i-���/�Y̵yXeCp�
�j� e*�:A�SZ�xy>���J�aWL�9��Y?���[X�W4�]��d�v6ұPzQ��J
���w�-��S� ݮ����$�%-�k!iZ�r�˕5@�;\��N+`�u�x�WE"W�o�O�vЈu��f��=�}e�g�fJܲ�-@�χ�V�O��'ۆx[ڶ+<������D>�/u�D��[��u��*]@�9֕y_��JWz���5�lu�c��5��=.9{�}�e�����ɽ�N�y�d�~h�đ4�,mF��p�~���v)��$P��lt�lT>�I"	���IQ_���$L�a����1]��W^���������0��O�?>^ ���w��������~������P����7w��/�+i� l�H�4��K/`�1/�ATP��/��:¹�E�I0rF*�����L��Pt��.����9OU%//_�����8�o#7A�� �h�lT�Y$$���H����$�H�	r�7H�a�mD���uȔ��Lʓ����`r��	;��D&ܮ&`��״*{l���<�	�*�0�/Km��ZvhX��
��Z"��3�K�# ˔#���*"�]�1vܶ9аUBX\'!��$`H�!3� �/���	�6 L�B"F�AMo���nI�Ka�fڀ�N��L}�X��SGC��2�T��QR�uʹh����4r��ŘJ��%���a�:�^�O��ipx%r�u� 	��_���O��`���#1�:`�92Z�k���%0dfB���3\���l"Q��_�I�1���̯`]��^F�&0�i�����,���SN]&� ��\���� l��n�Qi��P$�q
R̆�T0�+��kB�<�\Iñq���d�m�H��1�N��=Y�� /6�|�:�"4�^���}�m	y^�x�y��vfSϕ��l�)�5^�]�0���5>�|��\�~E�/�k���;"���[o�����te����)��ɽ�a8ȿ�wvv�oon���tV���|~Mҗ�l�%��i��H���:x��P/V���7����^{�u��._����Y,�.�P�bH���A�P�T����(�2-��MT��1a��1	34�������    IDAT�U.dD�`���R�6s<�B�Q�0�id�7ob�z@#��&"&���������Q�M�G�˩��4c����&Z�[��JN��@6�C'��5,5��"%�JBp�1ӡ5�%�#'�h:MRt�2v� c�F��� X@��F#s1��u�+���o�JzV�L�i'!�Zթ$b�j[�0��#�cv�2��Q�7�+*B�$b�UHB���q�`�Ev���f@;�UC�1��k�5ȧ�6���S�DY\��<q>���2�h<�e�;����cT�h[��-�55z��%�I��J8��	�������lD�SqtL�#��=oR6��,�d���v���,�V���\�m�f�����dB$+�C�o���'���qG	���{:�l�T�׆=����� [�=����k�,�Z�)[�,�)�N��-�Y�l�MoCJS�7M���'�k_>�O��}�
ܿ{�33�{�҅�l�>�q��g��w��f��Cj��R!��@T�H��n���i"����s��#�Z.Ґ��s�vQ���$��RĬ��DE�=%���bm����7��uK����^?��M�7ĸ�h!����I ��N�B i?ǈγ�P��_�_{��\xf�\$�8J���S+��"ӈ	��
cО��Kc�a���8k˄�9�z�;!��pf�SOMT�Ԫ:tv���kӯ�m�N�Fw��j@T0�FY�Ό�x ���\ �v��q���@ 2`'.�7Ҙ�DYR������e6��u9i�1����댦�f�s6�,������D����}�3��$5훔�È^���gk����j���Ѡ>E>�7��U�/I����:Hⴐ7O���F�	����86j{P�i��8ⷄ�qZ�83��1��F��K�����!̚8Oʀ�:BBHJ��Y�<R����hێ��;�f�rn�u�	�Neulk�����<�2�ca��L�l�F���f���s4����7�ŀ����vdğf�]���mN�`j���=#�Z�q*`1�}�Gt����aBmq��[*�񵍵_y�����ڇx_�������G�\��I^�$����Mꎁ�ј�~,3�g�I�����
y��=I���sBRĞ��Nnʒ���i?a�7Q��\؏)�T�.�yհ��71���.ۦ%S[�1�ɍ�e4D�c���$:�U"CX�*
Zg���f����ذ5}�lT�M/��¬ͤ��o�5B���F/�����pSS���F�Q���66`�5C�;#V;Q��$�ZCTC�5T������٫�RԤ��>0u..Ĥ��29[��uN"ӷl�3�<e��L�����FR��ݳ�=Y#$����&}�=��mۄ�+c�X�0��#0%�%n�(�C"`��I�����E_X�#Ge�����	���p\�~��+�@�	ةؔ^~��9��d?g_��]�=ȁ���@wx�������LF��K%��X(��T	dR��4��P�s�D�Yj0���kl#~{�ς�u�Q�]7ܖM#g�Nv}��Z��{ǈ���+a�Y�%Y����IS#���#[�}�l)���>& ���(�t��-;/<te�S?m ������׾�����C�����[M8ԙ��縬p*�NFGw��Ŧ�����F��ϔ3!�i�`��Me۬SUr%��C2�MO"E$H֠ns0�x5M����q%�~J}�S�r]�+PT_?�����h%���$ꈥVLs�7�����f�Q@���j*V�o�r$�����T\���ޓ5�h�e����YS�uF
AL��)�ͤD%�v��T[r$�LE�_�+Xo�t�g�A$��O�]H�T+�U�H�%Ӭ4��?U�zM=K�^��H�4Q�!Id�1�r��j��NG'j���gӁY�x�.wH�.�y�M���JO�DZz����*$B�IP�W-`��1���v��&,�<�Q^'�8�1���t4�JL7�!��X4���\o��G���ᜲ�K��Md���O��c�7{�d%"3����b�6�,�xdץ=/�h�Fx���N/N+�S���Me�ulr�e^#]WpSޡ3��O������:Y��-{�-��}&7#됱�F��5��j��ө�	3[Jf��-!U�����&SY:L�8KD5��\Of��͞'SN��t��f��'>!ٻ�3 �W�JDa���W7���3�o|�߸��WW1�b��+���,`�x�7��P>��5%�!)�M�l�ѻ���Iհ]g�91 ���u�ry��4���5YT i�P�!�Jҩ&E�1h�r]��$ulHD���� �Ɯ-5|_ZHt�-A��i|�Pf��k���Í�k$d+
p��?�D�B^�	~Ph������e�J;��$�Sc���߲}hl݋��v�7�"�S.OSx$Mi}��$ړԶ�e����(��!�3k��g����i�:�6b9^�Z�4ǩf�#MJ:L���Y��)�jR��h��ؑ��~���gE[�Q������Z�<��,!D2� �R��~ �H]��P��N]�>\3�J�@�FĚH���<M]$i��.:A<����v�.H$�ߝ���ڙ,�M5�u ΍![q�J×�S�����S�#��Ҷ���Y0�v#J��3tp�Kf�h��}*iz�)2�+Ζp*�&�����~^��� �e%�˙�g)�'��06�d�L�i�IIN�E��Y��!��;�VIU`{�IYs��^�1�L�p���W`?~�:2!K������r�0F��c�=6�H���X��f���r~���K����Ǉ>����~�_l\��7Wέ`�e@��3�+RQ��o�x��E��\�ڰ.�ӣ.���� R���YZO����c#����z�+#5ڈ�b��L_kQ-��3�D�'{����C��ٔ��4Ȝ�-�^�&'[4;�YȶL$6�c�[�'ӎa&M�cY�r�I�2�O�T�[S�����K4;�oU���A�K�b�(G�����M� J���8E��4~�{��]aK�T6�l3a��qL"�o�X�iϥ��I���.h�#����޶+���%eʠ��;5�B3�QJ�J�ʺ6�l��Ð�d��Ah��k��dM�M�+���^��y�dQ`�r���3牘'�kDAd�L��n�l���q
;K��_J�m]�,h��*���F;b� {V�(f��~1
�EU����G�0�%���Y�&�d�����W���F�F��\�q�����ҵ�j�a�zŤP#N���5��ͦ�J���k`�-����(�k�% �|�Ym�J���)�I����̧d�l)���Q��t{���^<��P��h����z��ʟ}��6�^�Of��sДToxI��N�48V�LQ�>�v�$#!?u�t�%�3�7��8�˦�.�'	�*�gH=&�f���P��h�ɍ9�4O_Z��e��7��M��D�7�%Ai�8�۾n�_Ҽ"��!�<x�|H�e{W3iz_�
�V#qRX�D��ک��m�u)#&�(��F�B�~��ɘ�q�����:��͂#��Cj�&�GkF�A�AH2j�iŤXa�Ɏ��Sj�ڞe{oD�`�W:7�5%����k۶C�K�w$`cj��9�R�z�:=) !Αi��\��H%=?i��f<	T4b�N�f��T"\S��Կm��X��zڵy�YWڤ`�lq.��*���R3&�| dr����$$�kE9!.�r����V9+[_�smׂ�?i%�t�e��ʕ^�O���c3�"S��ڸu��P���n�T����排�a��	�tx��A�$��>$�.�J%V�+���2k��4�u-��~�ӟ�n�{)�#}�a���v6�6W^XX��)�ۉ��i?�������g��ڕ+��h`��~�$�]�Ŋ��&��燀���mh������Mkk)d+K���f��xT˳QL�N���)X����51�8�f��q*WR���ʦ$O7غ�z�޿��������9�Ƶ�5�b�i~aXA�J�d�L�xl�`�=0�  �ϊ��!� ����c<���{%�Qe�R��
O$�F5kC�IqR�Xڰ�W\���k��ĵ�P&YbU�9��;v,�I�~x�r���f�0L�e����ә����=��:1�k���H������w&���FƲ�35ahY��,��Fj��t5J��%ub�87�,{O�P�hi��c>�,��w	G�mϻɤ���j9 ��[�E#o��B�3��m�co��1�33���i�Օ�m�����|�0�Je��~Aցo�q�D��r���hLĴY��4�e����{x�'�79Q��F��-����f]^^��~��O��>��?��?^>���R	G'mT���)sMys&x���鞍x� �1��W��l��E�z�b�Ǟ�x)�H�DZ7�g�����{
�m_g�Eu�M�Y1�G��, eA��g��_��H�4	�A�k_�흎|����/+7(�*#�0�V&}-�3l�!�T��>u<�L�_�WY�bЄ�;i7�z�IK�a�Ξ�1���,�*@�@*���4�B�K����@�6k˴��qPD��L�M��f��H4/����^#�w���A ;���}�����e�O֏�/��0�v_��σ֨��c�7Ձ���W�V�1�P^���(����:Hh��5	I-���̽�k�5�'UG[?�R��k��<��6��-�0bV�Rfܴ�nF�f���U�@�3�A��1��r���ۢ�lץ���7�o���#8q��4�̈6����O|��!$���95�=��Lc���pa��ɕ���~R�����x���������Q�%����6p���5�%�6D�j�jo^E�E%�UB�x3���S�xٞ�~�7Ӂ��p&����)�̮
c���Ѓ����|��߬�9�3g��مi����'d��7�9��"l��D.��	�k�D.�Q'��r�ykȳ��$�"�[��Y���EL�D"�2��j�X��Sg?o�~�N�ݟS��]�Q9%#��ޤ�ib�SQ�"F*P�ȁ�
��h��m�h�N��T�6�>tjZx~�����r���A�@����̡͌���e/�=&�A�8i�k��x�.x��}"�7fxƺas3� ��p�0�2��HW���%N��&?#��@�kLA��5� uc��u���z�>k�]{M�U-�ĉ��l�G��X�C�l�q�0���ߦ���ص)���4�{��jΗ�2��K���4iu�5"�nmm��#�X�4�>�(q�r�c���3�^^^~���O��>�����/�������!��K+�F�/�ۈ�Z-�
�ʨ1ⵂ�x�8���� ���(�	2d%x-�9kl�^����8U�<{a��C�5 F2�� �y֐d�G�Y�y
3?`��F�A�ekV�0gA7�؈9�|�%�S`>fL��������|�V����t#�o�uL���uD�'�&3�G�D�lvĉ0}�V�?+�8v��N�Q�2�K���8{��5f��f�׏�$�$9��:�%��7�Pgd-�$24�f�G���R(�Tt8NQ��A�$��X�Mm#Ks0�}b��R�C#X[+��t��"MM]ײP��&�t��Ǫ���$�T��0'9[b�|��k���jń@05<I���ʒ�=f{��T$��8M/�*��}ٖ�mP�ҁp(ޣן�mD���T����T���3#e�c��تR���L=vL1dQ�9��M�e�q��HM�}9���>��l�5^��O����?�I����z��ދ���++������|N�F���r���ͦ���bgX::�SسF�����$LM�;��Y��t��xYW� �<(�|P���2�g�;��V��e_���cl��>h����������8��SY��n�Ԙ��� �R�c�w:�������ˤ�&�ղ�M�R�Q��l��=����w)Qh��k����`������;&�'�1�h<�����흶׊�|%����$��o�i��ڰ�lȐ��҆9
�T�rl��JX2U���^���xd�Y�Щ@:I��<�e��(��G6�y��ۿ��'�;RD��`)3��`��i�]�WR��5u��,H��S%�[ވ�����𘎺h�ۛ�f�x���6
�rލs&��c��U2t|�(��b����a������J�+�ޒl#o�v���ܭ�u���3#br`h��rޱD�T�ⵡ�ۻ2,j�~����Ύ��jF��lU�|t[�q�;7=��kkk�~�'�sz�}�Ņ�������6�W$R啘"�
��\�i&xE�� �ޔ�G�3-Vِ`h�8�X��(=�dX��m�9���W���bF�=��zT� xf���X�X�wt����9�������')@��-pL"�SD�A�����X������_6�2��6R]�qː�u��t6ړAL�O{�4�ۤ�h������CM���J��,��?kF�e�2������@���<F���o-xg{B�{��N�IA۶3[��^[��tU�?�+f'�d5�e���LfN�95���b:�^PL����Y�]09��}f�����;+cUǜ=���?e���8�L�[�]6 <mJ��ȷ��<����Y�2���N�@�s�]����y��i���� � U��6�i=�	����iK��Q��u�-��}��"�}����##������4�:8_*bzzF��A%|�8I
�L�Q�A_��ҥK��e7�N�p��N�ccc�������=�>������˿z���R��M0!<�+�s�6�'�f�" ���Lb����Q��$��M�̺�76O8ӣT��|��٦A�1�eRM6�*<�S,c<M��M�e���f�����.;'�o��ٖ��gSj��$�U�HI��^DLۊu#��Z���'o����X��R& ���˴m;|"i��q6j?����g���4�a�-���P�CTČ���M����; Y����e[@?��v��̡=��5PQ�")MF�v�E�;�~v��u�t���p[b�|��D�<�.dJ�g�Т�����$d�Fq���Mۖ�1�L�qP��k��v߳�r��v-Fq(u}�#כ�3��wM��g��Q�"�&�#��IYD��<O�� ��n� ���шT��Beqƥ�>qJ��+'5�>��汓��v�O��mI]�$���@"�*�{,�e���a�m�	mEy�cq~���6�O���n�BA���0�;�u��(��m\����I�F�^g��9�muuKKKB��m-��>굊��g�ko���?z� ����=�~��翾v�򗎻�1����E#`h����^'����4z%�ں�ވjP�b�����b�X�q}�A�L/��I��F 3� %iB;���yL�P���Y�6��5ʧ������k�o�D �L!D����r\c֔��'�@ȺO&x�����̀rkܬÐ?;�����&��M���G���d�5��%�5 nARR�&�;K���ma����-��5]��4c��&r~\6��w��@��D�q��Ԏ�F2�x��6��p����?�VM�Umg[�d�M�Ħ�-��v4���o��\�H����y�L�S:���,Y�=�reE��(߳b���HFY�S$7��$JK�X,([:�����H?},���}�"%�)!�q��:
�
癣�>�o�&�4'S:ъL���O�71;����}��%�#\+�'@>���J�����8�0{{������|q4!�Y�_�S������k�9�fp��8�]�N����L3a�/|�i<��'������f"_�x������(}�w�2��A	����R*��_��;?���~��C��|�{�Z�v�)���K�x��:�q��x�Nd#^+�A�e*FR-ƨ��;1�d��K�*	Y-�I�z��g��Ƈ7�����l��Yi?{�dAj�IiV�J3�.�Y-�,����^@Kǂ����e-#�`I,�vd[�<��ٿ��l$v�������M��uex�Ti&ҵ_W%�q9v�5֡��5:n�    IDAT���Q��=�-�� ��ڪ����s�x�q�&�<�T�Q��5B������"*�f��ݙ�J������O֖e�f3���E���]�5>v|d(�e~F�D@ʞS� �u��]����pc2+ڨ��^Չ��)��u$YS$�HM�Hwg�B���������# ͈sȩ_�hLL�Dx�b��u�l�.�U��P
MH-���ܢ�o�G�܎0
�3MT�.�2�W���Qo����������*�Y��ts9ь�9��}�D�R	�à�Z�l&�5d��5�Rǥm	#������[9n��̔���ӹ`�J���3��: ~���� o��U�1O	]��w�1�����xa5S@�Xȡy��M��������{Wz^g���s�97Bw��9�lf��(K��G���z���r���*��S3;S���뤱d�eQY"%&�Q$��sD#�ܜ��y/n7��n�_���.4�{�������<�9���/��>������gڻ���I�,^��\��+&�����Jn����\Qjۢ�j�F��*��t�"^P��L���vF�U��aJ�y�n���#��������i5���{����m�v~���h�ߙyV3^�UU��o��R�R���M�d��5g�j�i���m�RQJ]UU��
�V����Y�z�ێMB�����_I��~>T_��f�V\1S�fT���s��}zQ�����fW�>���/���.T3�j ��������kQk��T[ժ��TK��C���ۢ�*5_�Ū��j֯(`���T2pY�mE�
vx!�Za5���rH=tۦ�Zk��h�N���Vk�MŪi^��=�(Н�S����ܕ�6U
����\���U�Xe��X��~  &ϩf��	d�V�ʸɪP��5oG�b����yrog�iP2)Loғ/�1[͊S}��u�T�L^g ]�+Z"T�)�H�+�(�F�E�]Ơ����Ӎ�M�ڠ'�Ia��Ȋo�xʋ۞j	�zeW2r?�z��i+A��k۽�"���"��Lb�քս���F���f�+�ݽo�d2�~�Q�x�o����v8���W�f�����*��!�HO���?��
���u��ܥ��ڻ�J�+�f�/��ITD���ޝ5���m�i��Z5���yQ�mG��*�ꨐ��ϒM�H%��搈sg�l�A\ʝu�����J}e��o;��!����k{d���F��I3�<�V[�v�p���A*}}£U���3ם_����ɪ�y�����?�Y+tc�'`G�Z���l�Yx+5ӊ��үx�}���
5]Vn�6�JT�Tܹ+��s�m���촺~����
*sWw���#��_�w�Y��iQ��v��*u���L����'�����g�6���dNj-���P{)�Kjի��a�Ϫ�U�r����.  塚��@,|keĄU�LV W�.���s�4����Hڈ������Ug��T�bd�2x������O+��{�_�6+ RT$˫�T�C�`M���5�ߓ�����e�D�,�+�v�\	Rt䳅� IեKbE���-�����ihM�<��|)Si
MVR%-Yޢ��JN�2a��Z�)U��sZ�9D�ԹSLF�3�(H�c:
J�"-D�-p0�m�&�Ţ�ڐ�@A|���H�V��&Ke���H$���ו��<&���J��L�+�JEv184�3�<˾��dr��Ǫ��L^�Ū�f��
{#�B>-ٺ�|:I)����ݟ�E��qz�=s������"��&S��xŗ�^��'H[X/7|.�!��P(�(d2�2iҩ�X�D<J&���0� w�f ��=�;_9�u���J-�z�*�wY�Y�����:�[�O�l�j��z��%�:���ȣRC���U����r����^���ݧ��*x�c'��3s�v����{�����L���j=U*S5��(S՜�{S]����듬�p�dTfy/��Q����E0*�R}��X����m�7�b@PqT�햑��U�B�V2S��ۥ�*e/aDe4Fx� [��˴+�W�j�Q���2��ba��X���x�0���&�*W�2�X@B�X2O�2��"���7��_��/V��{uR�⥽N��Q���H�mA�2�������*��{,��,�*&���^:X�R�C�����x;��\>��������Xk]��^�גL�_@����U9A���w��L&��2�ER�$y�h�tV=e}I}�$�=�9�l%2�����k��eF+�P�P(F.-���->�YɼM�l1�Nl}�R.�t�LF䋀3����l����ڎ����rb�ۈ��LLL��j����Q���{������KL��+-K>[�xe_d3��:o��8N߮]�!��8�(fW	�Ԅ�lN�rH���L&�V�R�Q��l2N.�~ax��O���/z�z�}���K]}}���2^�^�j���%J�I��u��f�+C귝bd�KR�$b1R��h�T<��eD`�L����m*��ZV�A��J�3˽��(��̝U����
����^��[�O��T��?gkW�)ܾ>��Td��S���F�
����I���*pU�^�y���a��W�|d8}Uxv?�Tc� ���fJ���c��_KdEE��Im���ު��
NTG��� ��c��Y��n���T�V��۞szO�^�TJ�m��0ʽ��v���"v̀d9T�تx���W2�
�^�6�K֣ƽɞ�v:�w8Ȉ;�[)��sw���'�R ���lSf���g���V�Ѳ֨��e���%=���բH��2�G�>�
X$,d��(�|�re�Z�tU@��r�+nO*2l��U�@������jKLu�J�&�q�s5��ڥ^158WZvtZ���M@E �QL��'�El�
�7��ˇ��o�6Uj�i�:�<nJ�<��d.�Fl��6�֦��9��a��w�3ۙ_�3�fla���L}W?Z������[���K���RE
Y=�`+e�4�w�w�X�{���,�d�\:ECM ��@��b�� o����G]>���8zk�����r�����on�Z�C=�T�n�G#7�]��W_����ӊ�\�`Ǡ��'�bh�n;ʁ�UЪ9��u���'�����=+�q^��J&#�N�d���~Q �e}܇x�;s�r׮�a�vwR͒��G��+�Z����@f��*�э5^{�e�B�(qEY@H%��-�m7�J=W���e����nX�v��/kՋUfu�WjʊFV�8�J4)Y�v#�d"y9ԶM
���j_�������P����u����$�����x�]���%W�Z8���� ���VT���ZU�1����VN���2Y'�D�(M�UڍT.�$چ���;%n��m�CT:"U�R.�YI�W�0�87Ȓ�Ц%iӒ�(J�o��E�}��)���g�n*"@���a{"M�����=�xT��* Vۤ�\�=���le�+5���� ��E�&Rǉ�R�j�jƩ�6��ݏ*&0jm峴�+��k��%��7�O�P�!���6��d(��DFZ��R�"�����LAoQY[�,�I=�D�x8M&Y�XZZ�	Y��B�l"B6���V�\1���e*���wj�d1������ۭ �l6�ڡdSf�E��ttt��zp�޾}���~��ъ��lR �v�)�3l���ϖh����؀�����B��g���]X�T�����:�~��N������i�r�QƇzp8-���fj~���Y��8%s���,>�m��<^.ݙcn#��|�pV������J]K'�����Dh=9=[k)L�ʘ8t�8#��𵿧ߢ�N^Y���U�����o�����j����խ5���>���466���/����*�X��Ǐ�^�@MP���|p��g�q��)V���	S"���Re{�)���������+&DX�{=��^IB^���%	�3R�Ƶ~�*����v=��
���u��ܥ�W�[[�H����_�d����r���f	�No�`+�"�T�o<�5�W�ن�F���V�	U�ڮ���0�Lhre�Yq�*S2ŦŬ�a2Yd<�:r��� �E�h0Q���*KF�V֖:CEQ].fT֛ՙ(���rR�j���L"��(AAtv
�#jT��Ѡ%�I�����p.$��g�N��dґ+f0�*��B���k;Ӻ��-՚	�T��y�-�X\r؛�&��Dg�Ld)�E�Ӧ'��b2�0uʐD@Ȣ5P�y6�UԢ�܂ ���Ii�l6��$E]Zf�SC��T���j�l�Q O����S�HTb!����@��R�V��j��E+ڢ]^K&�%Z�Q������I���BM1��K�s����Z��.�U�+��lUԦXK6*�j=1�z�YF�	��S�]8���6	4� S�[�w��z^��)�T��ׁ�n����2�4[k��Y�ep��,���z�<"�S��d�zq�m��iL�b�խu
�"F����Z3E�/f6CInߜav����CM����nʙ2��3�g)Ɗh��F47���Ћ�eR�S�S[�m&,F^���!*W���H+Z�Dkw'�-�\vj���|�2�u�tw�(������ݸq�W_�1��>�]���yp�&'Ǚ�� �p��u��A�--����1v�:S7�[��\����c7��=8H__���"�.��\:��a&�`��y�_}���<�����b���V4�}�|����Kl����#%|�v�u�iho�#O}�/�+Lܞ������G�au�R�x��	���=ƿ�ÿ@��d��Ώ���Nʅ"{����?��_�-��,���w�f��~.;{�#�����/�Ne�������t*c�K.����x��wX]^��"��d|`:�B৞z�'������5Чd����V�be�*Et����������c�EHD��F��9���/��>������W����$�y�j�khP@�jWJU`llTe����p�i2Wzs)���_cn~�ň�b��Ia�j[¯�h[�aB�Eg�\��s�L�\S@'��HL$����N[�n�;�4F�z̉pB#�	�EQ:R� ��DAG���h0�`׉�R�#-���ԫ0�͛)�����hC)`��5��!��]^ ]Z���@��Z}�t>��f�l{W�������^�P�Dj<�P�D,���V��=�D2Gy}��*��.��jB.�T�I"���ɣ��it8tZ��ߙL*C��@:�#���wZ(b4	���2���H���-nesG�L^�'�ʐ�执u��g�yk�e%�)���DWsDV�������O�(��E�4��<��&VR����RӔ�Eo"�I��+YRKk+��Zf#~� \�p$��;{���P�Tq2�F�ܺy]emK���O�WJe��[�8�LL�i��ߋۢ�e5b�Ǧ3DV#,NΠMg�	�X��� ӳ3������tv���`����D��RؚL{؛�=2E��1&'C\_G_߅����Ǐ;Ѐ��a��<[3l.�����׸�[47u����ݥ�5Ej}�&����:�Z�$L���ק5i�����L[g�z���;w�����*T�˫(M�xGGG�ɫ/+��`�+�VOW7��{�����\:{���N��$�=���:�x�ɇ8��w�{��X���9j,�nC�<��O�/|���yF���;z��H]����ӿ�y����Yؘ��62����o�[�ű�<��o���l�͈���/b�5�������>�Y����ܹ2��G?�w��&i|�]5�����Y��ϾBri�����^�=����jj����?����?!����o��:q���@o7u\�~���2��+K<t�
��N�
`n߼�[o�ə�giaQiYT���-ҩP�d:Óy��{���&ն��X['���[Q1r_��*ZQBK`���8|��ݝ�l��"����e�_��?�����˗[������dZ�d�����A��W;��E4�j�zb�n(d��7��ƍk�B[8-&��$.�Q	3�㻤�P�ҲyL-6�^��E8AqL��`"U��j�M@�6�P���S���'��cv��k��ۻ�ʀ��3�����O���6�K��ų�cYt%e�462���SLR�D(%C�L��J�����>��|Z����::�Z��}
H$P��V�L	(�FU恵���0��Z����k�z�}6WVU�%5p�|DY�/"����L��LkC@e���t<Ehe���E<z=u��6,z#�d�P2A\�Ϩ��릭%@�8�R�R.�f"�r6���G�Ã9����*��\Ͳ�Q��lKC����ɬ�d�����&�c��U��F�hR�+�ь�������-���͎�`V���rŞPS����Է6c�z�˥"�յu�� �����Ү2^9��l`��^��O9��{�`�})mlm-�*�[�X'��R�$9~h�I��e���geq��z���Y4��� .m�:����.\��2���e� ��T��j��S�P���4K��%Wq4�t�q7;p��К-\�3��r�SW�)��pt����inÂ������05��#Ѝ�ӌ�`��^��\=������Mj��V3��G~���YΟ;�p�RZ�ik�oh����a��^�zCݣ�6�Se�RC�l���S|��_�.��j�5����������������	����\��k�����?��SS\|�=LI�WG	�X4j�����}�ܺ}��GF8w�6���:�R��~��\>�>3�SX�v�f�y����k�{l?go\���ym?>5�sp?����G��$��.������c���kċ�Mףזx��r�g�������s�m:j�؅q3Y��'?�˯��Zh�G�|�wϼ�� X���Q�������T�X:�ɇ�b�U��fgme���g>����yńH�V޴0w:-���?�ɓ'1�̊ڗn��e���S�͎�fU��f8��tES[[�G?�b�Dx�n��=���_��}���s.����RD�	jk��D}2�/�N311��.^�([d�NX\����
�^�p�|2��b�9��j0�t�U��Z-�9Ra��.��L(*H�'�=���l^	V�>'n�	�Q�(g��n��,��-Ej��Եy�zdKY2�ˑ,�f���-��ɛ���~J+�����r[)��,N_;:����b4�E1�Bfc]6N�a�g�b�iJ�QK<�$�Kc��=���f,N;�WQ�Rk�v횢=z�$�--
�E`��'�v�*����*k�=Jؓ��Uf���B��@C�K��JSЃY�~�(8amv��w�����&�y�~?K[���Y6�i%����h�u��Ǖ�rx�[!�=k�{��]�O�ci.��R��Z45�d�Nt���i��-DX��"�����liDc�`�;�d�֧ak���5^�M��475��31y���@2����#�67bv��hnW����;�w��a����'���gg�T���oW�q{[������z��Z��� �\���t��RΧ84����/���F1�"����% �NÇ����٫J��+�����l�b7�����KgY�Z&e�Qt�ih��d��觡��W�8Mh��Zd��a�i�����|�~�4���,Ĉ%�4w����O��lr��?�˫c��yt�8-u5���>���޺�k/����P����`��^\^G���������L�)����𫌷��K��>��������M�Y����g�ڗ��p� ��5�;���q�r�x��J���-\Y#��%�%���>���m�ߺBS[�3c*�u��h4v�w����|x�H1IJ�$���`��7�u1������x���}�	k�lzz�{s�ɛL�,����0�jT��t�#�8F�� �8Ů�zUJ� ^2ڙ�IB�M���J�>p �߃�i!�
E�u�6�x\�C'Q��yU��V�_|���~��J �/
#��]������1%`�[��(��z�R>#���5�N�
����|Wã�>�$	����;�������/z�z�����{�FB�8�t��`�R�J =x" ���R��IW�+}�҃f.��s_e~~�s�^Zb'    IDAT�cu~���z��pXL*�~E�����
�$>���S&��!s�-�:�)0�hh���0a-�T f��u�P��ÍɝG��,3Y~vw���	�>��Z
zZ��|����"�(����^�:b{�1��X"�>�6�F��B�݌Il��I��')�QO��Z;Z1:-�����@C�W��؉�x}>U�[ 4@˿7o�_���NM�q��g3�ͨuFc ��`��h���^��k7t��m,�Y�_d��4��FK�d��d�粳^cfs�0y��M�h�b5���B+���l��e��l�l����L���"���d���%ow���U�dd5���:��Vg+Z[Zs �ťXB��B��n�����H.������ȍ�W�55��G[OV���j�m��L�L�����#��u��J�߯2��Q>����w���s��Y>șS(ejo��Ez�8yb?+<��#�y��^��Kcd��]�kj�r�ɦ�|�>���������xT���䧯���@��!�z�e�Vp5{��L��O��@K��]�������5���L���'I;�Ե��h?����ؚS.8�S�<D^����B���G�����'h!���ӯ�_����ַ��׉Q��Z#���;�������^�)��`���V��.����f^�rIѤ��_��TZ����|�ُb0����ߠ���B*��n�\�z�	����W$��i����hsY���[�dj~��O4#X���2a5�k�M�Y��1YE4��_��FO��Hɔg)bz�̝93�1|��Ɂ����𳾸���&�M3锇���������e�PX�"3Ozsb���z\&���%؊�S�k�mm�o��.;���M4�֝�lE�N<���/���t<�+���O^~I9O�\��0j�;W2��w�w9��LLNO�TW��"��6���b�Q�aJ�*ӏ�v���W����奱C���� ����=�w��Ů���ͭ0�\�@M�jё��пҷ�����1>��Ѣ6��t�a�"�x�,.�3q�&w����Bc0��nQ�j��SJ歕5³K�6�x1Qg�᧌�n"�ϳ��ʒ�ii��g7�1�qX��5%��L'�(�4�;���̸kumz�<޺��D̈�kx����,b�"�����B9��V��f2� Z�}f]|md���4�N.}��C.5�Pܼ��N����>ں۱�lX]��UܺuKedG����N�չ��_���q�զ����m����R��j\Vv��R��6p�LR9V&g	M-�K�iq�ir����1H�2���)d0��t46�X�������f~k�5B��t4�lub�iH�r,,f�Z�w'���4�%R֣��ɤ�,Oo�0�Br-���Ec�A�)M9�eӤF�e�H�ݥ����]�j�hM �"o���:���{��r*�M2���f��zWZ:�{����Z�wn�dzz�����V�?O�)�4��?�#���o���٧�d��z�8~h[�K|��>�ų�|�2�u�\z�mڭ6�$�HDU�/���Z�����4=]�kl����؃\}�uƖg���ù������k�����+o�Q�;�^��+34�<H�������Gy�?"��&�231���l
r��1Zj�����&���}��������#*���w��֢�.T�I����;�>�N��s���)�`x�,V�PI\�U��}��jV::�����x���ܘ4%���Ec��]K�߭4w�\!�C�������3`.��{�D���,/`�א*f���&h�P�� ���1���\*��F�7��ހ˓��ұ�0���Ɯ�+�t���փ����&�c���u�?�u��)9И8�Z����ר+'�$6h����W%�f#�b���9�n��:�V��ۮhwa�n��a#�����ر*�jUp���7���?��2���	(a�d�ʀC�W �G�G�u�+�V"�T��V]��j�"⓲���\p����ch`P��s3��G���w3�e��������{��Ŏ�]#�pT��)e%�IT�⪲������+��R���-�\�7^{�۷o��������nk�>��e5`��	�HGV7�ϭ�Y٢��d��M,�U�%�J��d#�!�-1����:�B�ER�,�ufS�]%�{}�w����X�f�B	&�2�?c,���=�.�BZgGc���]��1�Dq�������x�M��Ő��zsj������F��v�B�x&�v;b�����A�F��"m*�CN���#���Sk)��Lƹ~�*/���?8C0১���ׯ*AQ:�C|�[��(�<px�C���{���&�f��$�!��ɣ��[��Ե�z�,�,0�<��iS£���0�7��xT�t%�ND�֠��c��uY�oIg���0�qq�L�����?A�ldfeS��q�~$��l��#����u�Z'�p��ӯSc�c�Eh	��jlbue���5���_�h�c0h��V�zbj��(�E���	��VI�S>|��]�N�X�U���o~_}ܵ���)��_���������>�͋g�mo��[2�(O=�$wo���{�8�=���{���6���́G����+��96z���N�V����!&F�sky���C����v`q�48�45p��]�V4�]+��x��c�ݵ���t4�p��u�I�lF�x}�A���6���Ϋ�!V����b���Rb���z��{���4���#GG0[��l�z�x��W���xd�AZ[۱Y+t�{ff�x�ͷx��7�E�*c������h�s��u�v��#�w�T��b.S�s��٫�	�����qq�58�E�~�d���E�7y����>3��&A��T1���"s��&7���8jJ�-�8�f�bi�N'����Nʋf�!�f/e)����V���2M~K����n9�jT�D�i�ۘ%>q��r�]��Mu�W�UyH�5����2�������z�1�,ح&6�b���eu]��F�;�t5�:�$�1�|�M^~�E}��k��3같%	�(]ǧ?�i���'Jj�J+e�ta(zߪ��P�RC�yE�|aٷ�ө�V&��'��s�����C�\�r���g�F(L8S��*�U㳴��1����e�f� ��1G�%(2~��.�#��r��Yz;�i�1�����ZL�i2�8��-RK[��x��qF/]@擄cQV�a��iU�z���bq�"���̆��I�Q�h�n�wo��:F����0�+I�ͥ�M[�\��J"KAk'+�4�Nb!Jj%C��I��26��&M���K8!t�%?���� ��}��L,�"	c��T3���?��O?���g����bU !Ѱ�C=vBe���ϥ����[������OߠW�����/}I)��f(����Ml��Q~�7?���<�=�}��w��ǳ$W��3�FWm=�?ű#�z�-f槩ijR��>�.�����mW��x��i
�"K��C���"�)�)�vm��KinG���f��_#����L*Y��7�RJ�)��d����p��m����V�s���ե ��!�����t"��'UC����/�pڔH������!t-=�M��	F���Z��ڣ��P͒)�9}J�|�������௭�����O��wy�ͷy�#Op��)F����$�Mp���N��>�����+�m���Ţ�P��F�����K��w039Ξ�]��Ft�"�F/3K\_���� ��3x�G�LM���A���eFǓ\_,p3bĿ�Iw������]`el���,��Wp���#��4��rs�0�V�k��h%e�r���e+��T��������X�8�v���
x����OSSM��K�W�����R5K_������j-��L��N�[	�;�Ge��|�:�S������ޚÚ(2\׊Mt��5n�-66��Lz�:��
8�	̦"�R���*����F��ԡw�0��1;�l$�\��re�Ϊ���㌧
��.5�+�3g��"��]�bl:6f�*7����[bo�����^���j�f7�NGY^���sq�G�����j6�r;�e���V�6h��T}�R��W��L"�믿��fa
������E,v����Z��FFT+��ȋfC�WG�Ŭ|�vg�k��A i�:�9��` /����ɑ}{�4͎	�Z�[������~�j}SӞh4N4�dffFeR2�+T�xHˏ�GU#��j�2eH6��f���s��֘�}���v\���{�_�x��|�o��&�Ë������a�9�(��{��6���Vװx��E���C�a�N��F�J�Y���f�X�b�ޑ���i
��E]�r7�g<R��ӟ������/c��3=��̝r�����|��������oP�(��Mݤ�RV ��~����÷��uj�~�^�N"�"P�l5p�c|�ӟ�埼FkG;�+k�)�E�l>�ꅮ��N��[�op��Y>��{���3�������+_�*��<��Č��ч���ϟ��w��ُ>������^����xs�{�nnfi~�c��$��ƙ3��54ą��9y�tVz���g�`��7x�����/10\KCw�fl� �����M]#o�X�ݹ��_}v��7_~��FC���J��O�&7n�������7���:�lN��T[C*g߾������V@���[��0zQ{�����!����~z���,���^���-�_�\}m6��Z���O*������3O>���4�A{�To���BW(qὋu6����P_��2�p�{و�Y\�$�ɫ��ޮF�.Qgq׸X�opgm��.���B�@-�Z���Y��V�s�6��wR�{$骣hvc7��lf�u��sI��
�:�6^S�������o�����q�O��@�fֲ����ֲ݆�v��b4���R%���M�'��}y��aU�ڝ*㕬mmy��~�"���7��D�!�&��Q�S�H�����GpX5��E�f=V���w�]*���~�K+��6�q���-�������}C�[X�l�2�l��D�+[����P3��nG�C�j����$�f��0|��X�dQ��l!�b����2��^j:�ҭe0�1S�_'5}[x�#�n�ҩw0i����ɤ��-Oh��ēc�z(���A��iW�O)-�,3��C��(�J�i���o��/��CU9p`�/|�����bV�����*��+T���q��'Է�J2��]z���o�~j|�\J\���4�gϐ o�W�>��{�ƭ[��M��pLm���Y%��XS42�S|��=���5�� ��!����"�wX�����K�ߋŬ���<�ѧy�{���k�v��׿���>�8q��qzF�p��Y�g�pjXmq��0���ؼr����en.L�0����(C���u|���i�n'��n�l��ur~r�O~GKHcGw��3q{g����{�>��G��g�ǩ	��e���<2�����<��Q:��8����g�?��O	��������g��ݬnn�?4���&�.]"��� e��C���V������Q�~p���i���Pu�`P�b���!��������ԳOs���飫���ȯ}�\9u�7�
CM]���+�k��m���:N<���i��y��G��O^偣G��A٩����7�r��\-nb�10܀�΂�g��	p��m�bz�K���am��br������dm.B���ٙ�棄S(��}��z�ish)�M��\���Q��6��=�������W�__K��z�A��lf&gfT� �{��Qzz����Zׯ]Qt�_��_)@1h�*1Z�j�d�=��1�I!��r���ƹkh#)�s�4P/���<v��p2��ܚ���ɱo�.��F[�6�1ƶ�i�ؚmt���+�s�(a%����u�/��.�b�?J��L��¦�_�s����G&G%}#���L|�6,��^fw���AG1��n1�X��Z#�RO�� =�}h�E�.F�A���N(U�(z�`�(�@������c��;=9Nx+���5�J9�����'��rQ�֊�p�Ƅ*����ǈLN���#`�4c��D�f�:��;2H:��6��M��R��x���'��>�D83�ú��i`=V��d��sN��L�f2Q U,c5Y�.��:�Jj�D�O�	�Mn�39�]��򋷱��8�^�pK�.�UT��禐������������}h�:e�"%�T�j^X^bp�������ŧ4
��;o��O~�����ad}�f�*�<��kj(�*5]�⧻?�Z��R��d���K��ϫ�!����AS,J�4;4�'������+��\�������Uv615SqXI%T=�n2S��gM%������څYE��r�۷�1?9��i��Ə^WR���|�;�nq�g�8�6�K��<}�&vwu��n���>«k,���������릥%@<�D�]�Q�N�2��A^y�e��6�w�P����hee)̭��y7/��Mϑ���l�a®�\�6�����]���jkGp��Y��88���ȩ}��~�1��������2�k�������7���3<x��/�a��A�j"�{G����̙�j�B��2�hmoS��x<�]Z\�?���P[�Z�dx�o��o`���ۿ�K~�ӟ��^��h��B1��#�٘_��O���~^}�[�ml�k0)��Cȕ2���?�kW?��w��R��im���:66׸9}��_Kޚd�P3��ۂ��fll��u�L���bj�E���m#��\g}!�!�"�ar�%Q��3��l�|�����9|䨷9p[L�)�ڛ�u��w����6Z�z�[��L�ddiuU� ��ttt)��d�j_��������3ɤڃB�J�F!�S�]1ŉ��iZЖ��=KF�Lߜ <��#�gOM5-�bN��$rfVØ4�"��}�[��Ee�'�Dx��bg��]�Z�x2�MiJf�H�y��*g�,��q�~��-H�����Y�0ui��B�g&g7�R��ƈ�P��5Gz���'z;�s��a���	�C�m�c�уt����'��xQ�S�p��(��G{��0��UZ��e����+<���<�أ�� �>3��+�$M9���A>�ɧ�GVHEV���T�3wg��;s4Y�|��Cl�ck�uh�L,-BOcw'{G�ID�)���4d5fb!n�Ct��mo��$�:6������).LZ*��If2�+밚�$V7Y]%2]�6��w���<Z��x�Gg),�E�2��:7}/k�SJT��:I%#lƄIs�7<�[�W�2G��ɥҊ�_Y]�kW/{���=+m>B5�:��W^���>��k�928Ag��D�"r{�^���Ӵ k+ ,@m2���`���J����{��w�������.��V�F��~|�3�3.�n���O�����ؘ���:�+y�w�x-�f�)@"J_���r`6�X]�����v.+f�87����Gt}���I�n��\��UC�b�`���ݢ��P$ʞO�o~���V�^�b���:��w�f	��pq�2�=�.J�<um�l���>f:f�'�A�#g��Ե���&�i��p�ݻ8�ĳ&�v��-t�\z��|��/|��7բͦ������Tf{��i=�������v���T�Rf�J}7�H�����Ȉ�I`"�~��I[ǥs������5�j��nɍ��s�:��8Jlk�=�Zh��`�h�;��ci� �/��8s�=���Y�r9u�4%���&%>�f}�-�Vr�0;tj.���q{m���c�}P4�)�����]�sm��~,��I[\�zr%3�l�$ٜJc��br�'Vt �n����-t˓8�˴Y��YD�S���-�(�p�x�?����.4&6��!ul���AJ@�'����Ue��do�LN(����/+ǟ��ֽY�6�Y�,���G[J1��A�ߌ���m�(�]�e��������8�Y,�&m�\��r,KJ�;L��A_
�Ӥ0�5$5E�B�L'7�����Pzg��6F�Xb#��+�|0�f��G��O2/Q0�q,D��L^� ��Ŷ?    IDAT#�~�����_�c1��>=zOz��ޏ%�fmaM)�٤!���Y��X��'����d2��I�r��7n��ƓO=��PZ9��^���W_~��}���ڳ���O_��L
H�RʰoO���ǉl.�
��6?}I�����ǩ3����D�'ILMP�!��3��l�Kۚ��C>��U�.�g*���h�����z)�Wq:�p�Ml&����̨�k������J<e�8ImDY����x�Z�>��>�i���c��D�),�R^��k��e��H`��q�mĢ�
x�N+���Է�`qK�׬�U�w��es+DϮ>��2ӂ����$���ҏ�η���R��D2�>�'"�x*��?�y�6�B��Lc5��U�w�PT�]	�$���<_(���{�%�׳����v��jkk�����^ևxO]�r����?��U���^��N2esM�ż;��٧ư���g�(�bܸx�A��f�f�1dZUI��ė��n&)�G�q��(�Ő���������V#�tu�(U���T6tM���2Q����@�P#5�N2�-,N�[9nLŹ����Z	�zѲgM#���'71glL��P���CB+f���u2swi5Av~����RMf�1l.+�D�H2��ί���wu)�zOe�:��J��Լ�#G����U1J/�I�⌎���ď^x��ϣn�h"��A2%I��5^�"�M�ߎݪ�*���w�_#=��=Q����l&`�^�4Y]���9�ż�p��!Z&���ΐ�qc�-O�i�`h��y�{��)O�Xbe5���,�u�l��ڇI[�$Ż�`dnr�ŉ��|��$��h�-��h��8�;8�+t�4:��3Y�F�Г#������wr��h�륨+c7��2T&�&���#O?�����M����ys��v�a�gz�'af�A  @� I��I��*Y�u��e���-��d�je��%Q\�@��0	�C��}s|s��睆�� `WuM�t�������;O8�9����e��>y�s�����.ϓw�M��d%����}�+-ee���Le�k��d@�����_�4�s�
�j^��F�c����(���[/�1B��ZҶ�q���n�p����hR�z_�����c��
����?��q�[P2p�}<��	�]�W�Q���^�D4����.�������ۯ�=�?~�8pa���P�4�.��o���y^���t�����{|�����e��3r�}I�T��?��������8:�goXڻ,k;XZ�¯�k�z5��b�6���[���OPd��r��!�Z�$+{�kTQ�]�Fqzy��@O��4t��6���8��y�>�E���
>y��O	h��H�_DK-�8����=nc��.zk��_�'�#�Ԡ�>���G� Wױ4��t6��v5֎���QcZ^��K+�]Z��O3^��X��Z�x,�?��+�\&.�x�uZm�ş�����<<���0�B�ʚ�����dA�!�Y�oi�\��M#�=`�u�6F��y$���K�/��GG�å����p���9^��޾sdb��Fhu�\v!�%����p,���S6$xnEF�G�UJ�,�λ8�x
����`�A7R�1��GmkrӅ\�c1?�� B]蚈 !*D� '8�<�rр��L\�^�c�[Ƕׁ>S��bcg
P�mDB�fK��m&���<sqia&�D��jc��1��}X`z�Mxr�Vd;����q�l� �^�,t��}4�j�.��:��f�&N/-���6ͦ���zm>A&�c����t��J^ā���g�}��_�F��W�C��28���6��Oϣ����e�
LU`�3�Ox��
A�y��IUE!�aj"ډ���t$������
t͇,�<���`��m���W��i=v�9������� �|���hK9؂3S���v� :
11�*��(q��rU@>^C����!��X(aժ0��'D<Oyܮ@��x냯bv�,��EƤR��N����M4[-|������g^�t�Q���?��������gp|p� -S��4���ܹ�Ss#�w��-e%Tw֑S����>��ݧUs��w�����nc�L=j��W�(

�|��_Ck���.2�����^�Z���+�x��p�C�bT��C�Y����h���_��w��*&������'Oao��x� hsX��!�9h����	�z��}|��k�&�WW�t���-4��B�|�L��fMjr�2����ci�|�(��Pu*U[�����������}��9��O���n��`�p�>g��#���7��}d�%�`}��^�wV�;	��OCm6Q��1�i�h��0=7��Ôm�����š��j���c8m�0��6 q��zb��3��Y��������:xz{�v���W����A6L�Ȑ���`�	��>Δ3��f��A���&5���2�,V�\���"Ԍ
�TR�y7���wa{>ٟ>���Y*��N�Z�G��ٟrv�n���Q1W���o���+Ҭ�s�S� EA.[���8�T������1~R��t����G��#���r��9��_d��r������E�v�Ǧ�D�"�ڌ���`�K	�����iӑ�#q��&C.:ԛjV�sqjBh��m�)�p�l9+�P�a)?� ������a�U����C/^���!@�:P�m��z����c���f1vڀ��CPbԚ>ݰqcWŪ����+p�4��p�Q�Y�~z��NQK�������A�߃���U��#Mȓ�V`��%���g�kM�������3��AJRt�Ǐ�!W(0�wbf��!�Ь3e�?��`Qtr;9��!a�&B������I�[���P���&�ͻ!��=C��>2}�fΠ�ZP��,��&�U+�E!r�<��?���T���H�Z��V�EnyK��A*�!��T��qg��OvDנͽ�W�'�`��{���cx[,-�A=��J[0��%H����Ptjx��,��9�>�H�N*y����5!�4|�;����2�*��jZ�6v�vx���oa��l�A����&~�0����xx�>�wv�!+\����,N������ 0'�(�&V�b��S+9|��w�����F�{t��t�����／��[p�{(dXI��fk�Ư���+�K��ރ ƨ��[�񏏺h�.a��_��j��GVP�=hb��zO^~�~
�M�^�"���oރR�»�����n�gA�B���H
Tq����&�M��u�n��q�ӻ�o�q�b�b�+)������?2��0W$b�*��
8�0�ׯ�GA�Q�D�H�܍q�y���[,Oz&?�|��$y�
	A�N��8Dyrc�Ed�	2����Z���~[���+�(/��+kU���Z�;�l�YS��C�x	V���*$QE��£k��&g^ES�"5� �}��]X���Vp*ob��a$�pF�e,����>�cX������:�@�Vz�$X�F�VΟ���%��J �O��Ii}�!��R�K����9|��ڗ�rn��!�����\�h�)�!ॲ�'7oa|r�ef	x������o�r|<;9�R(�.�s��/5�����J���B��������%sf��jh���.�6,	J�5���l�<hb��@����S#��a�51
q�����$874�كi;��RV�A����@�k�r��Ć�w�J!����v�Bш�so]@f$ �u9	�G��� 65L��>�� *~�#J�Z������u�>@'(�2�`[rV��c��=\���v ������Nm����4^z�F�Ē��HX�2ލ�M�f��^eV��<lO��T.%��W�����m�� ����tľ��r��%��_����4Q�a|����lrs�!�����z���&1`�;��E	����Η_����w�\J2�k�C�y-]���R��/x5c㠋�;.>9�@YxکW��&�y'�n��Q����ꕯ!_��g�}ԭ�A�n�޼�Ѥ�^~ú���?a_`ihu���}�y|�7~�疱w���.��j1���n3��/��̂�Q
���o��/�;��;��_�u|�ч�X]�!ьd�f���������[H�t�ȊRZj~���Gk(D޹|9���QES����m�8Z�7>���8M�+����Z���p����9Q����j�=��,�G��u�Ѱ��GA3�ܮ��ZE�a�ċ��E��a^!�B��}�	��X�����d��,�R�0���9��֛�;��gy���j�q��}�r���k�D@�j��8����������6MC��Θ;n���sgg���)�2�!��ȓM�=�� t�9l�T#��k����s��!c�A"��5�ץi� /O�|�@vT@��!�2�!�ٸ�.�:a�"�� "Y����u<����15��!�HZ`A:ZC�S����dr��3̟���G�����8�be2|�"<|����e�Z8���vШ�y����G�7Lj��)���S�����̒�˥f^]39�% &���)W+�u�S���{�����/��/�t����0;u>���>����/�O�}�/]R�*�:����?��c#��׎��{���<@�b��Û����h($"���}�*����E���.�[��+]$�q��ܺò��1�v����R_��u4�w�EL9B��c��)�UW&q�k����	�L�J��	�?�`�����a�4c�)��juq��#�+���/}��n]K>���6��>��Ky���q��v�ƙ����g���߆�+��{kD�bp}��Ro�uã##*�G�F��wn�Ư~���?����7&	��f�`���"~��_�ݧ���Bd��~��{���o����q�9� `�ZE�sY������8��x�	�v�ie�q#�g���_A���w R|l;���N%L��҅��j��h�����o5ѭ����%lE�Z����:Oo�dU��W�`�0���m&We��>��u�G
x��cnq�{��Ds�1��.�%�{��g'�:"��m�������������;���?B�V�
9��R>B�S#x�+�ar(�^���ލ��X�� e_ĵ�\�PPD���Z��&�����B�����œF���,ξ2�Y[��p�>.��˛}�ʋ�.��va�j@U�;ؿ�o�u���\q2���.��>�g7a�w���2�C5�JB--#�kU!�	���;l0���l�IR�d'w��-���q�G&	<c�!`����Cf4���ap` 5����G��b�J&b.�_ċ� �$�(@��ύp�t�O�0�e0K��`Z���mԭ.D)���F�I�Y�(�-����z
0��$�!�<�G�;�[�-�?���C+o�q3,��EԷ�xtkQ;���W�#��<j�D}��[��\c�X����J$`��v���n��2V^8���eP%���LO�w
�._���
hN��v��x��l�:g�T:�3���F0:1�4����<�S�c1���0I�̙3�K����ﰖ6U4S�����ڣ����^unj����H���9^�O�=�S|A�3�X��bv1�@��=pp��i���$��L	x��&�+��"=ƷP�_ǻo\�����S!x}� �q#r_{�u4���=ڇ!����n�(�9X�W��6z�
�^�3_�c��ǽ:�g�q���
��ށ�	�l�x���ޞ��xSo�
�CG��DR �>�~r�Ch������p ��.dI��>�X݁v������^XFج�pkCAϷQo7�rژ^���w�@i�̦	�&%�%�����ho~�:F����+�Pzc}?�����'7��w�C�Y���"��p�����g���_�.h4�`*G�O6qxw���[/���`}"�h	d����!����K_~]@��Ô�\��8¶�Dqq/�s�t�(;pE�5��D�dO&��<�v�!bY�&���UG}����oA�WP��p�B���w�.��&��8��lV��E�.�n5Q��Ћ�z�L�ϱM��	���b���[���7?���,t��%wG��������}LMN`{{�62 �?j����i�wv��J�?�����0;.�Ma�|�ɍ(� i:6Z-u����Y�@Vva*	9A=�c��Ķ�F��/N#3@θ������V��o�X�v�%�sC3EDA��ݻ�HH�y����a�d�*Z{6��=ƫSC�m�frE���=��V{�����{��H�t#����|��-L�N�L(:$�\�A�Ѩ3)퓏?���8vv� �?�"��m�0����˧pay��rUFA��=T7vp�hSz#��QEG>NG
ے��Z��0>:���U��KT�jb������(��&r�YD�7��k���:��*��s�����ITY;<����[���e��8)��n��3X�� �:&�o�:�Pд�ȗ�X8wS�\	��*x$�B�w"9H���Lg��On�rδ����
�����_A�T����R�T��UÞ��P`Oej�����{c{6;E]<����	>�v6������?ǰ���o�ʗ%�|����>[�T;>�$Q��zt��c0a�n�vV�f6�B��U�~������8�I���;hcH4p�p����"D���N��,�ͯ����BpZ��~Gv�;�se\��+�O
��g�� ����k��p�Lc��7�T��J�0� ��͇���H�f/|�0��O�\�֫ �~
���E�fǐKĎ�������[L����/bz~A�ݓ����HE�$1F7����L
$�������=�|�n<���J���`Ʃ�Q|��1PP! ��Wַ���#��,�L����a}(�������"7<�KWΡ�� x.W:��ݩ`�&q�._� �hC�V`G=�"�ۋ�/k0u�y-1A�yX��o��^m ?u�~}��D�B�h�=x; <ù�<��2��+8T�u�����7߹���IȚ��;*׻���A;;�x���`jr�K��N���4��� ����J[`�����P5",N���++)��E�D<�[_݆�����$
��2��|���z�^��3X85��������l��X��P>���S�
6
C찏Æ������)�.C����+���{!:Gml}��p�����y
�d��WJ,���cЪ��1�rf�33+��o�ڇ�T|���Q��/Aճ̄'�O>��S������;P`L���[��Ec�#�U�x���kT!`V���42� S#sr �۾�#���K���l��*�q�UIP.e1=5$�Hĳ��1v�{��	&�'����!f)䐰�i�֓6;ԑE���F�"l��mW��ք���<De�	}Iք��W�Vv!�>ی�g^'�R�v��*I)��e�M��P�LSミz��;ۜ`���u\,��~e��V�kk���{�˧�too��;���5����-f�C��@�"��	|� V3=��Se�4
��9�(ba~��C��k��ų/�͍m�x?�+p�ɓ[�b���88�`}c�v�7�G�ae�,�g�����Z��?��!��H��f�4Y�� T�Vqyi�]�ש�ˀ���z�uC�g��4�0m&��#��*�҅^��K��#Nh��j�Q�ɘ�3o\@qZ�Yn#�-��7���j��h�s�ae��J�T2{v��>⚊����
�|U�, �UC�����=�8;3r��!r�v�˥�.����3�[�g��n%)zX[��B�$I�ÑY����������S�iӜ �/�_���s��x�(eU��I���Q����G1&pvpf���w�,a�Y�^���p+���!���c���X�7��������(f���^���?�F��_�4Z�    IDAT�?r^n��ꩊ��=��z��.
S� �g�w���,4!���E�>��6�(�b��X�����&.bx���̃��)�,G�ǨVk,9:2�YY�E �7�?��������ν7
Xh�'�S����H	��
J	9=�.��]�����������4�n���� N��ZG�����9,.�C'yȌ�0��-l��X�41����I�f�]��Z�Ǉw�����  '@ؿM]@�(A�r�ժ��~g�F���D$��S�!�������`��V��& �}T���{���Fs���^������)@�13��
ԍ70�x�����B��*-��;ܧ䞸N*j=�$�O�KLf[�����0�&P�h숕!񜾃��m46�����\��m���\4�X�I�2[����r�Y�4�pZ�
2#d�L�fI�'h�:�p����C,N@�/��s��_�G�Ё���0$��P�`�D6:�w��k��yE�.�2��I0�&���-q2��Le`:�Xן>�,��d*�	��6�99��s��>����@Q����q��U���!�kΞK�rf��ǹ��5UG�DHF��G���340 CS����������W&''�?ǰ����'7��UQ�qxT����5������=�3�x����6(R��꼁	ӈ�@�Ce=�=8�C��"rj�{u$�*Z;U�vj��"V��tz(2B/�pԮ�@F��/BWbd��"D��N�ZUc:�^<����������d�=�F�.��0�4�3��z�����K�����)2�*�]x[1t�ӳ[���@�N���h�}�.L��s��H�mE�砨xwk~�ʕ+���a���i-I�������{��<�O�&: U�kU�Oy����(��سx޵����1��qa�4�z���*T�>g�4+{��%X��QYAh���j���Rg���V���4�=<�@�y��,��(�H>1��Ml>ރ�������E�l�sЅro���0���0VF>a�u� ��u�6�aP���W�Ʌ�>�LO�p���#t�=|���8� ���󱷳���������dH�̎e#N^]P�kx���,�H�^$gֽg;��� c��02��� G�j?����z��a�OMa����C�v�`��Į���J3�G!�}d�}G�Oo���~e�2���"|��>��t���W[��_A$!�� H*�a/ck�S�
^����0�<"��344�W�P�ᥗ_Dix��*�Q��\6�������TC��)�$���o��o�у��Ҡ���rq�K�RBA�����ɱA��J�,�f� c��S�*u��.�3yS9��JM�Vv�A�怐h�S���Ԏ�uxB �lB� ��,�"��i�#7�b�����CPG����P%[��Щ9P�e�� ��,�W��7�Я#��Q��160��J�,P�w�I�AL��M[: �^��n��Vr�/w�e�+Ut�ΟZ`����|�Ѹ�5	�4�*&��"��2�d+���X6TU�@�"6!V.�E�x�$j���ryt�����߸8I
#��/<����'7��򋒢���f�6�o�2�(�%��˗.��n0��>8�,�T[�0�S�2r:P#��L$V��<J t���5azΎN� 6��B��$qQ�ڨ�����K+�d$�Q��b�[óV60{�4���Ī�V���>n�G��!�^EP��o���S�bgm��5M�g��HC�W��F�f�} �J~/���[=��� f��9z���f7Ϝ����Q,}�D�"�=��c�t���f���Z}.=Q����|��13=�����u��)N�)855�ׯ]d�#��G!�Aek;���,�8��丆A��`VG7�� u�fZ1��_�
9q`��4�n����6F΍a��,Ԃ�l�N�O�ww,�ܓ�L]�S���!v��$���-<����vó/A5��rR�C�*�}��C�@.�PT��{hvk�.����Ayp ��A&�A��xأ�u�Ɨ�x�����J�l�o����#�����'&���cz1�
��'S+���x�+o +��	�J"�pc��}J����" �l�!�+6�\�¹�S0� 	��1z���vG�_(c�� 2�fـ������� ����KC<ǫ��ӛ�h�XF"�e�
���XՇ�@ja"����(�8K�U����j3�{vv�rfa���UʊIkzuC��l���g,NL&�?��?�/��q6ڧ$r9�*O�cB�xv��ˢ�/ #��|����w\G^V1hf��͗�8����\�Hm"��b8A�Yc��/=o@4��pj��!%tlw��Ɉ��W~`�����k;��Xt����PP$�r��0�$�)�jǐ�ź���XP,$�4��Y)�$�>�O�U��z�\�#U��Z^14]��F����I��t=�{�a�z�_� �:aQ��J��'���ioRrB���I��d��8�!��!�V�����[+� �ړ�ӏ/<�>~��|i�eU?��x�6� �y|t���WΡT*�ɳ�,($C襺�~��7^SC&�I��jA#wCfw�I��I�<1�qa�.�A�h�]T��ξ��|N�Ih!��vyk������s;]�V�A2"Ի6֏\�\��c��^AX����e���>��+�]=D��bf���yt"�_�N��P�D�k��� �����ad��D������`lvg/,chl���"c��zR`E�p�/E�T
��zC$�w��6��]�j�od}�R�.3��ry�ӆШ\}T���ud"�a�z-�b+�XĀ��,�p��ed�zhA�h8��<3|n�秠�c��nPG��[xXQ!��F�їMPx�n����P�k���K0�����@����&Z� 4qaj�8�)�d��� ��#h��7�z�e)c�񴘈.������^B�X�As)t���)������ƭ[7091�d���]"�?�v&��x�����݆�����6����Ș�eQ�Q ��q�j��J���Ps�\���A��
�Ѭ�v�k(M�1<���3�K:�����X�a+���@*MB"�UՄ&���a��q�8 97�cd�������-D�#Hv�,��P��5�+d��}�q��̪n"S(�Br:�F�122G�L��Z@kt��M������h�����w�A&L�$�y�2F>Ś��$H�:gp?<�Lr�B�;�<|X��� ���@�*��&b� ��	d�^(���z�@����0�"�a�b:D�B��)A�U�91i�?�V1`�;7��AՆ���;�^#���3�p&R^���0�2�r�Xb�z�|i_нm�)�*�c(4����z���ƙ�%�5]af3���dI�v	�5�z�"ʼ)HLB$$��M��8�yO>���^y�+�S���e�xW��syp���q���ԛ>� D���@��F�P���vvwy��qRf3����t{P�WWfqf2%��8BN�;!�z��#�V��ӋP�3���"Nt�.��mHyg/���WaH|��꾅�v�)a��$�V�!g:��"��.vkn�9��0�_@TGd�'
7��V�[���:�P\�-��ux�M��#�nSY�9r��s-����G?p�-籸|�4|ڧ�F	x�kޙ�Y�����X�U����Kܺq���(2�Z��,AL�����S�X���P�\�b̲~�jO���1.�G-�;�-xb�vr�����gQ���~��p��F��W9�<���Q���DM�Q�íg�5H#KЧЃ�DR�!�n���hw�0w�>� 2���%�Hz8^�R����OA#D�6��AP�Ԡ�t�)&YÓV�#���(L�N1�# ɰ�u�j�ɟ<zLIrf�@"�� ��L���j�!��h��Y�ʹ
&vW7�87D!�`P6$ ���B	M�B���0T��!3�K-dy��B�،�D��q�<�x􌴨5��h ɐ7���q^͡�_E�H��ؾ�d���fsh�C�X|�w�H��a�-,rP�}rJ�l�(�\d�$� �7(ۥ5���I��~F-"�"�9c�$H��T.h�Z!
d�8#РroB��T���v��G�Ţ VUDV��T�%��&���м����(��IN��	)L�x���ĄJ��$2M�+�B�B"3.g�q��Xć�*E�X79�l6�HiF��`Z���J�������Ĥ*|t��u�SDbL+)y��� ��K�T��KӒ����}0߿�������>�?���8"`A�*B*�g؃��ktp��\�t��~���x��������b��=^e�HȠ�����*�E`蠣����*0d)H��1��+�T���U�za�B�=��6� A�D���5{6r�a�O��L]iVa"Y�h�8a	��p�K7�A��j�#�eg_Z���A�p�k{m�U<9���P�_Fd��gk�]��`�
!̡�613w�T@�,��;܂ҫ��{������D>G�!�q�%f҇^�x��,t#�ϳ.2�'���a�W���aȏ����ǟ����<�A�<b8٥Ѫc�����,��H�Ȯ1��Rڇ�vaU�H���,��p|�ĲX�/?:�#��&�Ǡ�!�k�۬CPu����ȁ1^���8�,�-�ŵ�U[�rsnrBi�p��C�t8vۅ*� 
#�c�N��o0�@{P�����hC��0�<�0(�����7�0����
���GɌpI��  �y���/R�26>¬z� �0
N!F�U�* ����I�@tx]J�:����M�fdK�:}��A׶���]8������Eח�P
*�āj �S��zz^�fۇ�H���"�SQ�da(���w$���������@y�r{�"�����C��%��e���2QRX�L�\�X<C�1����y��?�`�2-���
}��p&1p�2A����(d�%��EO�,�$�tYa�X!��C{7�kx��м:�J*)��'�4���'��v��������<K�O��`R�K� ���I�p6�z��8ۥ�	
R�F�2�7ҿ��ʨtL`ȕ���H�^��x�����t��ؓk����PE�0y6��G�Xd���%�N����2p���#r�4�&u+b����D!**��0�����}���,Ħ�||�3�{�������7J�"*�=y�J��%���B?���e�F�ŤITF>�y�����8](a��N"�V0�� E|+�ӱ�=w30?<�U�B�VI�.eQ�^"�v(ʪmݒ�s3a�B5��� gM%v���b�8�F=BG���Afpn$�x�	�mX��*�!��ϡO��؇D�K�*�����s�,�Gdr@"�T�5rY��;�t�:��O��؎�e���+����lۅg[X}����ghU�|(��EjM=����y� �z(:FK�$��-vy�Id������F1�j"�؉"F�gѧ[S���A�p�=G�br>�ey���96Hp�uj��1�n�a�@.��SMt<"�P�������D��+��#f@�L�䠋nʰ��P�;���|h`zn�.Ï���d�4��f����7"�PA??�+�>i>|� ���}/���gA�ɱQ���~��3梬`ll
��a]ݬ� ����4�L��A�5�$�!&���f�GR��`dr\1�  ����b�ު�@����	
�l�Bu��
*��t��m Q �YD4����&����BF�3��'Hs�	�e>�I�z�iV�8����+��f�R�IkI�6K��>W�h����Y�ր9-��!����$"�Q��#pC렳 �,�|��E���/�}p1���R���޴�_��A|�[�����:x��_d�г����M�2�T�'$�S��uHN@>�����OT�(���!栆\�U���		?�M�����9.�D?�֏֗^�&�-&�4Q�l�>��KߔU�ѳ9�\�����ޞ����rO¬/«��y��?�Aqh�[�B	G�v��Ղ,�%�dm��H�d�N�3:��H�Y��N��d� �݃��M���Y�zFrB�	~�C��eS��XB��t=�7��+�kAQL�P�j|�T�M4}�"�F3(�)(��"A�bu���v�f ��Q��EAE�ւ�w�x
��\Bi�J�#v��B�Ն�nb �A)�a�!�䲬`E��<��˥��'H��A��c����4FF��*�	 �K�v��tߪ5Ғ�f�o[�"g�O#k���]�q��i@cXVjTBj<�`%z�3 Q���TQ���8<E�E�'���`B��2�B�$"$�tF�(8|��{H|n����\>%޾c�����d�@�*�,�p,RL
8k�e4L����N�Sy�v�������<�� �l�G,pbJ�~�C�,��t>�耢�
j|v'i	�֊��t�y��j����.YTF�AK�㙉Q�n��02�DI��ʔU����Z�/�|���1�6�O�I�R�����˔䡪�:�v	���D���l�aÐl�Ȥ(�[��`�sn�x��Ǳ��f����$�(`Mt��Rʺu��˛ĸ��bPy��~��Q0��(i�R�#��I�����!�<�BNX��){�}L}Lz��{4B(1�'���8.3s"
��Q:��<���3H�U�K�8MX��ց�)ʹ�1��I	y�>�Z�t��_�)��9C�I"e��'*�t��i��{�gK�?����Y%��@� 	�?��!�=��7E�t�릵�~:�����v�y���5�U5(i/QO�YJ_1>3�B�۲���~������>�������Կ��D��gХh[S#m2k���x��B�3�~�!IA���ZL��$�t��;����j�P��˖�k��[>fǧ���߃�hn�`�T��� ?g�!�q�H�jdsߎ2�e"D� �?1�YT!!
CY$2E��z��'¡)�l�n@1��QV82��,���tݐ�
!�}�3�9����������J�d�G͎f�9���C�G��*���Ф��^��Id�}f�T��IT�b��%M�AB��Ƴ(3q,> ،��0�J�?�~�
9�A�fn"�mSO��J�>k�BґhxD�#$�Y�!s��5��Hz���r�zi�����T�spE:�"L>eX
+�U����DvB�|�(|�;�Y:pR�TvԦ��x&\����IY	���9���u��D�#�(�s��0�{��p���4)�	�aB�?�Rr/ �*0��3��@}�Hd��,�Yfz��,���L.���vҽAٴ")�j%�^��,oȏ��&N88���k"��PDQ΢z}2��˓��z�a��hs!�ynPB- ��I��hN|cy�P��xn��&ϋ?/�Ҟ�D��BJ��\� Ŭ�N� ��)�� "�H&J�yʎjg�qVJ w�)�P5,��N^G
���K�����=��@��u�!���K��Ǥ�q�^����S�9Nx�Vfॠ�{�ϳ�P>�֘�)z?W:2D�J�4�!�2�Aj�:���Xj���8��齤s�A����O&K�����~9\8���++g~����������0>5�k��gay�m�iC�A�}�N�Գ�<��q�/"�8H\�,&�1�z�"r�hﳉ�CC�,c�<đou� �f��c����D��Y�)�4!D�1��	"�@DQ8H��،~�p谊���bR�	w��|�qyt��|�@싐c���*��*����11��E�ѥ����zF�K��nhUKg%�(���B,[��� �2I�#|S:.t�z�X��G�ЋE
b��1P�*�R�}0�x��$`/�(��:�(^�m�E�Pț�>��J�$��s�K�T��h"    IDAT�J��/NY�Y�ݥ��0�Đ���!�L�\�0D(�	A�����s�����D�:�t�$`�g@�d*NNX�,K$Ҝ#�8� ����i���'5$:�t�ϫҚ�r=���0�ўdc���D�D�s�Y���ɕ���0�)�����'"�YR��d���_�7)��{�Գ�D�/da�|MtEJ3�n����]����tĄO%x
�/N}ZQS���^G^�O.�g��'`��aa�ĉ�0UU����-#�ƃ��S�J��'D@���@�K���F���TJ�^*���P�%&H����Jp@��KA(�7��/��O��t����r4m70��k���Ā$�d�'���=
J�e=L�f�O���>e��3�$%���(4�J��2��`�΀�k� ��.����Ot��tJ|p:�4h���ꂦrO��݅Ӌ�:=���k�~�����@N��|�^���k��������������QJ�7HJz�H}��UV��#^�<t R(ț)��*&�Y�&��>|�CS�C�L���G=-�零jdeGt~Ea��S&��q MX��YG���@8$�%@lE�V#._jzq"�Am)DL�E�D%6�S:���C/"0����1%i\���#*eh��8j�CB�k"�PT�g��3�%P_���%�&2eU<�~O%}*KR����Ⓘ���s�>:��@Hx9;�RrL�C	*S/�rev"�����P��G�{c�����,V!q�$dl�������\�INUz�t�qFI�ZR�Q��~)��Ϙƾ�AM`�����=�����i[!��;��V5)�����P #�{���;�������#B�6�=��J�K	l�#%� ��"x� Iͤ����PEdI���в,d�E�{�3z�5���iI���~G)�Q������f�H�umD1�[�J���,���io��#Ylf2:kr���4]��r6���p_5ˡ��������s�3`� <����@@�c.��>���i�=�E�L��3��`H�to�����ZZ�*h� s�M��}Č��	���!ÀG}��Y,!E�~�#"Y���Q�����.�=�s{��f�_U�$V~K�9�p��x��I˛�tM��`����̜~.�{|��>/-Se�A��E��sH�����{�����&^	eҤt�Q�M��a:�-
,9�x
�f������s_4���G7n|'��gN��ns��"6*'��Û��f�f����)�2!�IW���."�Vb�xr�&gT4�O=3PIN��i솲O"�(�F�LY'������ȃ��<�J�qdF���	Ӳ���TZ�4��\N����dZM�HrV�B��F�����,"�OY���d&$�2��B�$��uB�ᒺ��`@�s �9%����( �/p�9#�9s�,G��1��	W
 d)E�E��T�׶�Y�L�BY�%��7U�yE��D�.����"�~R�UTM���	�(5�<_[@�f�Q�/��;�Ϊ�_���͙�I!����{��H�7B��!�@0�� 	%)�E��^�%tI=@z�>sz����{���q�&��ϐ�3�m��yֳ�z�q�EKd0�T��|�t�Kp%�!�����;x�H�b@&��d������K�QU\�CoOrE�x9��(#+r�A�N�ޒ�J�#C�h���
u�b�R�h�iȩ9�
�~�"u������p	TM�3[B��I�8�[�M���?�T-d(�1�� �2�}IaB"8���"_ �F&9b�����%���&�NiL&��i�(���3�$%e�\�`�RI�T���Y�l*ߪתP��@c�4G���%׵��4M�2;��=��0�` ��:�}fB9�u��sY��4���aV���ZRUm�`�VsiE``	Wl�ȫ�t�GB�m�Hf�����YA�ӚGG�k���I'C@&0���;x�<[Z�E��7�1�g�ϲձ�/L"C��{��Lp$���z�3�q,����T�L��h�7�!b�{2� �A�K%4&h�y���qφ���]��6��h[	�F~��t�>!%
�M�Y1ާ~�,����Dch4D�׊e_#��/XEkK��A�Ғ�3�ܠދU!'j��$����#S0�?n�4� ���B��d $���*���|�&�"��v�d���a��.\���@㌢�wJ�'�1u���Y!�X��+�r�W���nb4�'T�k� ʏ"��=QG0	y"dy�7P^2�1�T������ֻͬ��!�7}&�a$��Ӊ0
V�y4��Q-VU	GC�ׅ�*��iT	N�/6`,2am�E��d�-��=;_��b)kz�d�Ԝ��
J��r�50�X�W���'��J���VRT̪B` �q@��bJ�x�Y��X���f�D�%ț��׎�arA-4�/$�tv���d�o4d0o��<I��)1��u�!�˸�7žl�6_'�"a��
��Iٔ�5���5�v�uڤy}x|E�	P�(>ݣ�_��y������݅|6�vG���[$lE�	�? ���AG*;V����ua«@��$ј����*�w^7^禤&H;��t�4Ԥ"��1�<
�>v6���ZL�����6q=()bZ�����������$7�ZV�l � �i7���0z^&:���|jq�	�V˂�e���j�Zh�2��5s��i�Ov"�!���)��A3^�N�[C ��E�l�6�'�ǥ
AA;Ī��������Lq���Ʀ�PD*j����a6f_��!�����z���W���Ͻ��]���Y;���$����Ny�!q����bh�5��L�����'��'H�N�IРC��0V�U��emn�ME��4ԦC/S���6#�}B�V���a3^-�~"�̈́��ra���Hd�|�� �����M}k}�:*Ѝ�7f��p��/�.Ѡ�SC��9U��sH��P�����ʓh����ؾ�p}2���{������>���s�����D�P��nH�k�؟��U��n��/�)�U�i$R4�I�B�~æe����X���D ����8v����"JU�SY]��K�8�^���J��/�75n��
�jEw�!.uwtJ����W
L�C��
+�`R�ߥSyxш�K���}�YR�ѦZB7~{^���TȐ%,L�n��皠Z��ߗ�Q"��la�v�Ȥ ���χwֶU=Q&�6�������I���W;��l����-l��`��@�2��ϏP&5�٠S�*(��!ۛD�XP��=��[T\ߵvm�H�ɰ�y�L����	���U�Aғ�W��f��c��b>@u]dIj�L5=f��}K�k����h������_��Y�\[�-�'��|���"ׅ�GP����FISч�����ݙ|���-7n<�}��!�Gn�ˎϭg1�l���I�{�o��ք'��Ӈ#G��63N�Td�2(0w#�(m�R��)S����S�a�
�H�ƾG����O�r��*�g�dX�6�Ո�]P�we���6��⅕��{(	1��ڍGB���qS��<�Z�����H���P]T�E��1�����Kh�5�F����>�b�8��c�Z����1���Nf3�T���d�fϔ�.IG$��!^LgU��~�d z,j���D8�����T�OBY!���2��h�9�Px��z;��t�n�DĞ+Y��
��a꘷nS�쒎��k�T�tw����Sϛ��j6T���ߪHأ/��������U���i�=ڐeb{����6,�]����׀ �*��1�Q��k��3(��g�R%ct3
�e`*Gw}�|�Te3[<��m�Yز�]�り{n�~�?�z����l	��|�?"#��+��R.�iF�,� fOME�֚���D�V�jcXґ n�0���W�)�ګ���+�>WZ���X����3{��rAޭ�u�ݿ~v��o9W��f2IF�xB�{��Ň����فX4���'�I#�u&�U���lJ�Y���!4�<�1
�#G>ײ��&M��=��F���� 7�zǋ�dr�v��==�j����3��Y��LÅ_"�dٔ��3U^0l|RIt�����j��Cc�^�JWy���u�����$n����D< aТe��.&ʈy�ˑ�;��^PI������:�ڟ�*�6 ��t��Lū
@%Y	4�7�Tƪ��X������nL�^�m-ѣv#1/!H��d�ht �:�7N2
�X�h��98BV��l?�靿�&ߔ�&x�Z��j�v.wpS�8�T���K9�f��c���x�{�=Lw�|O�\��j�������$�rF|���5pp��o�/�p�0��EMf��uP���"ù g�=UXҫ��aٷ�:��{��Fz�Y�ٿg�oPˈK��J���j��l�������E\�Q�~��v\�4����\�͵��(e2rM#�k�*���V�շ_�G���%����g]���"�g�V0�����x���1��[���&���|��m����<�׺�hƆ���sš��E��'��ؤ�V��p�W���X���B�����Ai�e��3�D��dg'ƴCgg�>�����/������������{q�W��ҠA�-��'��l�\AC�NU�,IQ%y�]��v�C�M�0����y;�dn^-zp���,�X6�ka�u�[�����֮�~ᾅ��bc�������[�!z��칶"�C��i�i��uߑ͝��zM����ա�q�zb|��t\B��<�� �.�eL�ޜ;7�YR�D�/�=?��r�f�ΊW	�O[�:��l��Xh d�2 ����i[,긍��b&�0��RЛH���\?��0?��L�,��_������;wg�v)�1xh�/�c�ڵI7H�u���]p$a��3L���#�<���5	��������%SBt���h0�t׃���&rRM��g�]���ӷ�9"���HIL�,�,����Y������s��EbB�P�]�Lx虬��2������+P�[6�	� ��d��>�N��&j.���|�n�Z�#�Y֋2����5����T�&�pS�tuyl\k|��m���Z�!vI����=�z{����`b�猺y:�B�)m�9���rP�ڣn���\Ǝ°����#�`�����c�>���� �?�߆�[se�{��':�ۏ�s�=5e�O8n�>��D�Q���/���a�"Ӊ^�f̤������LF%}�I"\D빲OzO� k��o�rj���e��p��� ��u�թs�%�&�پ/7��],�ￎ,b��?������r3A�jx�Ap�j}c�t�<�,�����p����M>T���?�Vk~�ރ}V~Q/ʅ�`��4�jb
�e�;6�󦷭��J�6��^}��i�KM���\*I�^f  ��Lm�ֆo{��|L%x����0��k���q�;5���~s�M^/�fn�|f	5>v��������xj�tm�vcw0��![���+�!���Hj��|/W�9�N�}S���`�z���u �+K1���&qЙ_c��d�s?%�	zz&����;m<�� ��"֐��,\N��Ǆ�ui{4�}�ϵطQ"]�'Ϊ�B�<M�"w�&�2�Pcߏ$L%]��#A�I�L�f� �G���a��%!���T2c�,1�mo]{�e2����3�Zْ�b��$n6q�|�����OU�~>���P�UF�ɠF�Q!t��W7�D�曽>e��o����9�w�}wԧ�}�r]C�V ����!�-WQ�G3٢�X05�$�:�.�EJ��!�i�2i��u�.S��_$W��k�����n>�V����P�5^7����̆3��Q��k7qA���c��,L��w.Xl��Y1�`�?�97:e�f3T�M���#��(]+3n���1��������m>�NE�����E\�VpdU�M��۹ޥ�����J)����_�Q�2��O�t���ݤX5��ع
B��s]��XKGӟ���L��d~o[����[ �d56�l��/	e"Wuwk�t��Y����S|/�9�ٓM�t_�[�j�\��Wa�y3LZ���*��
�� �{�dK�I��d���.٨��ML����H�R�kL�|�5���Zϖ-.ڢ�$=<Q,�,f[I�w�/�/�CexT9(i%�clSd8�0	�񉼓!��_X��Bf�&������8%��~=�ʭ�#��^V��[����K�t��<��-'A���9@�\H�X��\oRߵnrF�&�[*!�%3ҳ\��Y�\S�|�-S��*Q)�P�p����I�81�'�y�����]=}h3�qc�:�y���agCŻΝ����������l���t�R�uuKB�P� {�6�����82�G�f�o�ty*|{:;�q657k�s�f D�!��l\������O�U��2m_��j�j{��r�鳦p�����#���أrP�	�%,Ʉ���2��!QO/`b�fs� ���]e��������;��Ʉ�`�&4�|����&��9G�������d��6��l��
$�4�7T%|��3�h\�A$d�^���Ti[�����l���
j�h�17L�
��p�&���wj�UM`������!+�V��[C֣��UR&.8�Ц�Um�k�H�rmU-R1/r�KHs�8=���{92���ud�$�Bl`�^�M�Hm�K��J��k.�EPbO٠��5Űǯg���DF��~au����	d��$*;Y%R��Ϧ��#c�����!�2�������nY�� Gm�<��Ke9g�H�~���s�`�*��*�&yn͸י��d��6�Z)�P��#G*�Z�c����Xۦ`�~��7�Z��?��@��C(�G_o��Ur���>3��S�{��w}�������7�4i_��;�;��.���#�oK�l�/QN�6��U0h(���2��^WW��M�-��"K ��Z�qt޺�b��9˹u�Ƭ�9�?t�pG����s��&��M�}w:T�uH$2����5О��B�p+��54�@{>kvo���8MŽ��j��m�����d���J��6�I&��"Az{��A@�����kd�lx(���j�8C�2�4��'�1�E����Qȝs?��&����9���I��A�ڬ����@~n�U��d����>:��uF�c�k������ԃ$�2��6�qR�ٱހ�Y7�$x�Ǫ���W�D�R�������<�F'���&���Î��V�(�$L����&c�l�{ǩ\,��e%.4�䈺�r9_��w�y��y��p�bH%i:�"|���e]���5֖�7oS��j��LxX=��˄����h��DI��]AWO�!����$�?��&��m�W�R)#T���;^�`�U}Kk\��im�����lqߡ�	/e����@���I�*�b�(� ЛM#�:�l�m���'�u���k��P���;�³/������ȑ�C�=�S���͘~
�&D�ª*a������̸ٿո7T���.�I��x��q���_�h4g[Wk�n!G�9�V,�\#h�_�め��lO�6��NK�
ͩ܂w�����UPF�J���aq+��{>��<w��X/G�֓��j�����y�B�����k+�~��nM��6�E�QK���{劙�c�H3�N{��Mў�aH��:LOn@j$��Ғ�"�u��:S��~�	8n�w/[
~5f��Kx�5e�B�<.��;��w�n��Ƚ�&c�(�f;�]=h��C��/9ā�!���jY#IB�4�,� ukWY��UJ��%�RW�V�䗱M�]���W2����i��(d�_��4%G��$�M���M�(�����|Yڌd�����?Ӯʮ�ɳ�Z!<�J2&�L�Mjt���Ll���Hʨ�Sh�Gј�3�NOo��D�����\�j-�]�rA��f(��o<vF��U+V�m�%0��!�I    IDAT��P*i�/v<�|�Q�W���ʕ�5ז��j���V��ߝ�%������`���$nWU�6
Y�\��<Z22���bJ(�L�p��VM2�*>����*(�5��'�o����ټ{v�x��+�?���O���R�z\SC#�.[�b���-�U9^������6o2��{A�#a�x�;�� Ñ��Ҋ���a�p�6	-���*+oq�T�a�OZ#����c��C��2 E@��g	Gv��|b����1k��,�S�sA��<��EP��f��H<����̸�j�n������h]�U+�q�L�^��n01����@���v��p*7*ycg��_����ف�r�X3k�G��]ܠ���(�Ta����=�E��Ų��E�7�h���c�:��4�'���k5��Rs��~f3�G=A��Q1p9ȕ���5^��01��ʆ����W!�� Y鬀�Z������J��1�pI���y]Hv�e�C�%Ų�r(� ���x\���Qߏ�Դfh��*��S�b�Ye5�����M�Hr�e=1{�!��P$�u�ϗP�T�J<�����f܂��6���z���>|�h�y���Gf���	w��1�`���I��I�b�]v��������t�5��oҏW���F3)-��!�/?�����9C��A\l��dLDxu��a�{���\&�!sߕ ���ikzgPz������9���`O�VP�ȆJ|�oϔW^��{��r�s!CW]�[m������f};*���ο��룿Z���-'N�ꫥ�Y�JBzBP�~r܌�<b��>A�le�A7��>͗��7w�T�Dz�r���Kx��K����>�$�3��9���g
�o�*Z�:����i�s�$�Q:� �<��T$�	MeO�!�>�`�+HPa���Ù>����b��a�~S�����t�Y�����%&Nw�dP�9��
H�<y���&Xn
�������ff�J#Y-�l�%'4�Zre�����$I�#�z{��H��a�2Y�������Š�@XKx�����E!�@���oA��� ���RX�����z^K��ަ�l���;�V�����'X��5刁��L�3����E�۷zז�k܄y)x�t�sdr9]kVI��X��4���]ύ�E��̗���bf_��P��oxŰfi�h�=î��H�N%I&d����j|m�q�L}l����9�50H����RE��R���WEK�ü��'�c��`Lk+���Ur�ph`e>���b^�0	J�v��4�0b�,+��V����Eᕗ_DK}���h(���M��XZ��(M��	��/?�/<��4R���HGl뇗bfu�f�=Md�xMW	��Z���P��O�d!>k�M���}=J��zV�`VنD`��%�����ʢ�����^ݜ���'ϻs��w}��?���+���/��2(��Dzm;�I��H3�{�q���u��rC�r���=�I<Zs�!Z�	�C�Y�_,O���;T�+)]b𐭜YTNgj�?S��NP~bݒ\E'���/r�tC�=.<�Ӷ0!�*���#��vR��L�����\��"
��|3���U䡂5}�:�ڊ�U�&�1��s_�y�1w
f���ש:����om�v��kH��q�+Fn�
h�9*v��p��B�ȠX%:6��>�V8�0"{�H�#�Vf���M�2N��������2���q�"�	7�I�j��G�5����UaH7��#����7�R������иa����KĐ)dMG�Z�=J�iq@:���&���n����d�O8����a@/�J�OU[8D�lJg�{1�!��A��P"S�(�5�p���:��lhđ�eL��m��S;_�+��u�`;g.�5����"Z�qd�)T["��|��7a�x�7aS<v�=(eS(�S"g1�eb�I�3Y��5���I��w����bْ�x��G��A"L���Xd,��"��u�1GI;�秞B#�l)2�h����l:��幺Y�J�-ܮ�ֱM�n����!|&92�=dJ�
1��������@�i��l1QGORZ�_F�����j:C-t��rщw޺��v6T��q��ӟ^kF`���6���#::��JYm��<{c��N/7��4�*+R�����-M�5^L�H\�Hl��?oԯ����'e�z2U�	\�"X�� �m��~�gT^�X�Z�Y(�P%+�\1�c�(��F�؜�ӇA�9��	>/�=��	��֒�ܦ�T,a��_d��sM
��I���|k�.��V7��럓\�)��"F�C،I��`h3eG�2�L�\�J&�bu��4P�4#9����j�N�1���ɭy�e3���GC�˶y`�n�X�����N��.�kW��������(��i���9_�{���Lk��㼚�0 �����9������L%�s���6p�S�vA�%f�
"� �c� �/!Qߠ*�h�exN������$���d�%ļ�8u�n-
Dָ� U[H2)V�\�d�ݱ{���,�}�1&n�)rq �a�K�#�Շ��݁�ja���i%�������ӹ���5搃6�!45�ɧM��eK���>�Ih���I�d�l=�X�͍�E<q�1X��k<���1��QA��B�y7�﯒b�xM��F��gfb�j���76�Q�����D x͍M�WȖ'R"�mU\��k�
[:6�V��m�Q����e���"�����؈�[||��[6�x��+���ޛ��"���]�������-[�(RȉD�#�LX�l��-(C��N!n��(K�U���?,������t,jz�
�5o-K��~oɮ�e�І�,ގU#��-�F�
G���u�%�l�c��z$���Vشs����i���#��c��Q�m��F��{�9�3<�ؚ��6>�������g
<<V�V�h��0�]6�F���?�\&A�h���p�nMEdz�ܰ9�V��p�2����9Ҏ���/�V5gaP�k�{�A�����#z&)���.1��"�@�d4.��k��57a��!JH,k�lT�����;���
v�o���C=vb�=���lK��1�"Q��~S��t�\�uq���k�R)d�z4��4��l�Um�ZA����`�KH�^qб�ǲ�s�d��r&�V>����	��'RUD �L�����R_3/�^r>F︩�ǽ���է���0����n6٣�A\.ѥ|����:M�q&��������8+V,�>�!-��G2��"���A9����d/N<�L�vw��������(����y�8�*����,��e�]��w�m�\M4�=-�D;��M]$�>�c��}���%a�K�BS�,�}�L.����}�X�ڦ�j�خ*5��U�,�D�E��������;o������w��ﾺs]*�f�;��O�!�C ���g�����	"���x+�sAM�BXMЪ"_*V�gp�D.j_�{SV_���&H������^�3X�����g9O�MW�*x
�5�.�#Tl&�0`�_ۋt�j����*��S6���-!�TYf�|�p?:�dl����(|s2����a|
f.�:�U\�U���ݦ�6b�5`�Ͽ��7��g�)ك�e���K�e?���0qr�%$��'�.-u����s�=2��ڈ����de�"S)u�5��A6����I��rUG?k�!����}�����������hh��T�����h��,�Jx���1a��5jT?뜁V�"�f�CUx]	�gJ���i�T�k�O�eNA�� *�L���ŗ�j��!҅~��b�����ڊÏ>;�+r������g���5��+הlJ�.X��u���ZK����`Pf@6S�$i#Z�����X�~���^��v� 1����-^�������Ȧ*d's���Boo���r�D���k�-���܄c�$�<�Ѓ���h�@�d��m:h���l?<�G�75a��Ëy���RI��ף��Ɏ��Q�Z#E0ka���k,���A�vX9�]�u@D��(�b�~�*��������$��L����:�a�����HBx9:�"����[v��['n��������77���}���>�y�I-VJe��c�%����t�c=�Yy��V5EP%{*�r���|E��DV}�8L5S3��L�z���.-3�D.3+5g3}kKX,�W0��{���d*����3 )�_|Oe��&�Աr�����1Ad쏕(�!�慐����	E��q�a�����Ѩ�kbR��X�d�|��u���T��)+@)hXVqm��ʵ.V�sf���U���.\S�� A�m>�z{�j�*ɻx�C��ѣ��܄L>�>Y�20��L_W
��L㥿���>����]2,�\��h�?:���d����6^g���+ U�����0x�4jQ���8Z�]'�QS��+ӎ����t]8��9<�ʴ��N=�����A3��U7�R!����Wl��6�x�8)�!�����k�Q�&���ց�eJň
������C�(�S���q�)�`��G��ِ�BO=�G|��p�T�Q๋���հޥ��I�ϣ��I��o���o�9k�A�6����H�B�\�s>2��,cu�}�9�B�p�	�d�����Y��Ň��x�Tu�Ɩ���f�B+�������8�3��dp��"�P�R�r:�f��Ke� �K�T�`���E]c��y����#��>�1��)�� �O�l"4��lz�.YeO�φ8
$:eI�#�L��b�u�vÞ��E�uϦ�Mi�E؛'�-�%��L�x_�m�⣀�%W2�fZ÷ݖ�9��I�}�1����kC��7�_�zsom�'�>z�Oh��E$�S��$k�ޭf��۔� �y���t��L��;Bj]dRʘ�o~���*@׻q� �RA37E��{�Ln<�/��!zp�p�(��Îa��=���Y��%{���Ƀ�ykݡ�#��Y �u����ve�H{U��(UCh˗q��a����b�sQDc8��6��,[�=�DH����{b�]wEeA.��濅��|���9�,�'7���c���E�ƣ�����s��>x(~r�)赓k� �����d�9l�0�k�,�B��������rU}���DX�UD��3Ͽ��;��|�ةE%��z����۠e�0����X."��C],.�*�b	���k�q�����W#ȍ��?}o��CXAǧI8��|V�0*8@��R���y��ԯ�A����u(���� �{�mjD�RB�҂HQ*�Ԟ�kA�[�F�됬����fD	Y�K�m���/1r�P445�l��T�hL���(���PHv�i���~��;m�B�!˶�p�U�p�G`��톞tRZ�b:�e_.�n5��ǐQ#0a�D�&�^Q}�E�����c�B;���=����V��94 ��_|����x� pٴ+k�â����]�>��8��8K-�'��v��+���ܻ�ڃac��%3��_"���"l��d2���g���o��N;M��yw�%s�l ��H��,�� �� ��Cw:�C�<R���;���%"1)ht�����Q;p�=�3�`L���-l&�ċA]�s��KU�i�I.�^F�x�hx�s��I�쩟=_㑭v���z2����;��C����P-�6ʏ:P�C%\���tM�쇗]�E�ĉ��e=��x�ㆿ��{㽵+?�}�I�'����>D
y�9 �Ъ����+�m咪>�yBN�_x̐X���
%$�9��n�4-�T�쿨b���m�KK��X0�ѹX�ʎi>�$�ea�t:cd5�H��9�%�%�qӹG�n�e ���r�ꞒJ�We�<�qt��h+�$����F�ӱ?Ş?�)֔H��HĂH�i�-W^�:/�~�$��g�����}�����>�@4�s{���ݽ�K/A$S0�dr�l_��|e�_�6�J��[o��D8�)]�L̐��z{~s�����q�AbĈ(����ēO<����g�:��������Fm��hX~Ȳ6�K�knĵW]�ƑCQ
��)N�P)��@2�G�r�R	M��Dģ.�T0&Q���*�G�7�/���/���"��R&�:��Pɛ�8�89~-S���d�f;�0r�0U_}��������ձ�{s�{��WQH��=��"��h��	�g���!cǀd�A�|�p~���n��ӓ���G#�����W^FC(�-'n���܈/�X��D?��p����_�@Ʉ}iՉ`�Q����f|���0���z�
�dm��a����!���ƣ��Q��on���&L@o:��׬Ė�n�)S�U��;��[n�?��1���b��C8��#��q������1c�u(��8�?F������{!���EL��&c�I[ �,���G��6�"���=�+%�~��x���q����#A+���bu�/�T.��')t��u��z�g�Đ�Fԅ|(���++W�X� �#>�	�._��/85s/�L=_^�8����T���1���]��-A�	5��/�v(�s�����Y�=&�NӬ$���`@R2�	$TqOp���)5�{��i.!͆5|H�C�� �+ ������FQ�4��>��c�<�ʋ��z��W�g1�W��I�_���ޚ�[����O�|��Sh���RAP(�Z�u�z�v����R�T�	��!�י,��!ES��O�Xf�"��ɇ���˱�	H�V�dJFJb\q����qc@Ǩ��HNMf�I $]�b�����p�N�56{L���$R�ۚ���N�c�1mp\h��e�P�M����������]�5��^��h$N;�4�Z�E#��3��z�5����:�쿟���7��ߞ|s�ގd��|��j'��c��gb�CR-�L��7�Z;�⋁DT�ߣw݋��6�!��T������,W����W_/�e3�Co�F)AT>d�E����[�Ka�ig�чB!DO>#6��s��4�9�XX�zV-Y�춻����}�w1t�P2������`��;o��v�^�C��5x�Gѱf�z��Ώ>�x3Y�L��_?�s�8O<��֬]��Æ��'c�Q#5��r��s0����-��\�b9N��/0l���O����=]���\�	n�e��gol���������o��#����셼��W_}�f܌m����6�xc���3x��Wqօa��A��S�H����H��0,�3� �ޅ�&�Lr% �2��&�v����E*է����p�5���ˮ�v;�B���_|��3g⌟M�n{L���F�����v�����Kx��g��S��9�#ڐ�Ͽ�y�ݎ_�p&n���V����^ ����A�_���0�[�_����;�Cx�2�}�Q��w`t��x�(�Ȓ F��0�d���gO~P#�9� �>7���W|�D�p^ȯ	g\��H����T�r0��ys� ӗ������B>��?{죳�[Ң��U��F�- x�n&�̵K�g��4��XL���j�;w9��,�"V�����{'�9����"^	I:__���$�)I��AǏ�W~�?⒩��ओ>�����)��x��N��֫����rY`��~���,�N�(+�}�/��le2Ԩ�1'�����1��M�/�`�.�ЕO#If*%*dj�=��W�`��?���	x4w�����h��$ey�2Z@^��o�i#��@�X���`�e����b^�K�㜱��z���� Ǿ$<28�I�^�'�����m;˻�������\��]t�q��SmƬ��#�s.6�bs��nJ^�U��c������E�ו�a�2�6ƍ�]�@,�3�>K���s�O�pɥS���5+W��;����Dt�`B>�d�h�d[����q�9��ǧM�N�TZ����c��    IDAT��|셱��zn�3�!	��-��Ie���Hӱ*���i��S=���Cp���z�_}�y�AL�f:�����_��{,&|W=?�=�f�ժ�YAR���/�G�eW_���L��YG�[m�9N�|*6�j=g7�p2ߘ�_sõ:���=�m��=������[݆�{�hG���Nf]r%v�~�sԡz��=�L�t�����y�?��_x��{0c�����ʫ/�Y�cΜ9��f� ��Ӯ��H�Ϝ�5t�J$P�N��O#�a�7���N9���>]�]Kנ�ˣ��?�|�>� ����V��K/�O�<r�{{Q%�_�`��o��g�3g� D�(�M�^1+����j��X�ч8�_����������c���Q�����ѵz-��r	���U�ն�-��E�����˯[o��N:�r
O͚��� �՜�"W� �b�B���#�h�v0�����]��p���Q-��PटJ 9�4Ƒ,��.;c�]w���nRo<���Jk2��فf浜�HTT�׵�8���Q�oH�L�Kus��LH�&�Fl�ʸ}��B��G"Q�RIDI$$c�2%� �o79��N��t2j�K�#��-+aʴ��"
!��j��-�Q�7"7�]�uߏ.:o�O<m�J0���ǆ��W�7^�i��x��6������r(��Ͼ�$�5ǐ���9�N��|W��_�֡�>�j*��6S��#ݧ�[�UQ��)�I���V$���q#b_���C.@���|��=BJV:�:��ݞ�+�I~����ƫ�D�>�l&���vU����5=��Z��շ�6P6��/Q6�Є��L�և��LV�w��쇽99V�YZ�"��$�0ٱ� �J"VE�Z��w��_|��)��u~�T}��p�嗉z���!�M?o�M7�
�.R����o�:3n��TC��W�Y��ڌH0�XH$+�y�1�M�:RIT(����k�QYۍ9�O�7E*�CG6	�?�Cgw�ߌ���Y�a舍�l���ӯ�q�������2�~(���?�!�fM>'��$��m[������(�28㲋9?�����N�����k�P��S��i���]tVt�#�h�{��½��_��ιs��Řz��2b#;V1"+����.��-6�GN>/��2���G0o�<�U7&���7��+�<��;��x�����<�7ވU�"u�/�WO1j�磝����<b2\���Kx�����;bD��kjR�!�ڷ�~��ē�8]�N??�,L�|��~{,^�uM���Zӆ;���[f�(צ�L�7+W�@"^���(��`U�j\4{Bu1���k<r�ø��_�e�P���\x��>}:�l�=�!�F[6}���ՙ�a��v����TħO�^{5�օ�8�JAnh��Ę�*H���Ҥm���&N����F�`�������~�����b�u�K��E��b��?��k_�Պ�lT�9t��ns9U�s)c ݗB8L�zH�,����=b�z�tc�Lg����R��%-H�x榑�gm�0��h��$���lo?ɧ%�H�.g�@(�N_�M6ƣ���㋿�0$���ק����I��u����̓�� ��-��o���t�1�
[&��A��IqF�Z+f��
�Y�cbfX}JD�Q�o�����%!ߏ �%�y��8�/G__
mmm�Ց��	�� �7rm
�*F���Y�ܺz{��?�����TbAAg�
t�l1��"�nhĎ����o�=�]3f��W^���G��V�Uc�޾r%��Q�c� J�F��\��������^�z�6Ǒ���>,_���#G�Ĕ�X��
���(����e�*�}έ���1}��XZJcYo���+�h��zc����d�j�}�y(�CX��ɫ��͊��,�;�|��>mԢ
���g�8�4��9~c���cQD���E�	.�u�}���蟟!�Wo>�h��;λ�O9Cw�}�8HM��E�G�<�V����PLe���/0t�(�=�r�畧��i�~�Ą1��1A�d���=�Z�}��6D��щ���g|��b$�Y9&M�):�PD7��ps�^����?�|"��^���˘;or������1�z��l�I8���������Ϝ��Dk:�1��	sgݢ�m��K���/�N��:
�4��"x��1�e0�>�0tp�uw�V�x����;n�]�U>�O�S/�cƏWR���|��r9�}�{'�`άE�J�F��H]=
�/�ɧO���߉!#�c��`�ܹ������}3���.�~���N��s�^��F6�g��C�u�<���?p�eS1��C�)�A�W}a�KU�D5��ɧh �=�oEK��`������>�$���UQ{8h��Ƃ:�`���X�\~�!�deo�5Y�U�U�V�����ܤ~nG[;*D���\�9i9���ժ�S�7���>�m[-��|!+oI��[� �\��W3TleZ����G����%��M8V�Щ�@�.�L�˿!��������e}�%�纡���;��k/l��\4�;���C2YD��`�lңyǑ��*���0*�簗�8�-I2�M�B�8Y��%��y����P�1�k4������i7��)��i?%t������P��y�f�I��� '�*�$a���պr�,�����2�0�J���F�����e��w�EYbU(�ݮ�[y8���Z�s���ϸ�QaMWb�:�Y���y'֬^�h4,��cF���_ś/������1�Ƣ�R@)`���8�`l��<�U��P���އB2�K/�X����梔�������kP������P���`-��u&m�5<�P,�hG%B�\����7��|ם{�̹��-�a?�P��C�Z�8�H?���C���H��p#�}�M\:}��z+%t���ы�SN��S/F�6�ʛw�)ga��1����2]���CH�=ě��^;�W{�������"��t���'����E�c�L�2{6��ӓ�P���~�W�r�J�鉧0q��0�ι���w��>|����x�ч��_�ǝwމbcT�tr���pu�E�q��p�٧b������ᶻ��R�Y9���K>����p鴫���AO�L/�1�5�oo��8~r��
�������*x�o���o�=��A͸h�%�}�=q�q�k�]��p�_}�����~,��\9�
<��?�fk�C+�_�iӧ��W���#�{�M�{�=�a�Mj�T�*�4���7����}�!R'p��t�OO����}q��/��t�/�I]�xÔe������a?Đ��qô��Ic+��┳�P-#�"��[�X[�FM���fߢk(�������DoG����k���x)�a5�!��6�6!� ݗ��R#H>�����k������f�7mX�f��ۧ
Ŝ1��kژ�*�ݿe�a/�̩�&�ӎڔo��^���Ő
y���x❷�����c�נ�Bf}>��͹����[F��nړwߋa�<��,��^�&�9�	���ֲ��l�d]p��L�[aP��X*9�W�\��Ҝ�SC�
fb(�L#4#��������5x'� j��ѣ�{�9�pmV��zFR��8vB���R��-�﮲����ޯ�!p�5{������\
b�?�M&��~|:�eA��^�+������V[��=�bA쌕��D)������7p��P��еj-�q.��d�a�>������0玡��Q/��@��c.2흸�+P�"=��0k�-����ixd�f
i�&�q͕Ӱ�{b�@O!�<=�@!�ŠP���Y��D����&ٍR��hT���n����,�F�F�Kp˵׉�:n�$�v����c���b�//�OO�	6�m�fR���[���.��|&�M:!��r�<���<�����⩨5RU�>]���_����DDc�6i��=��?(����iW�ʛnPu���gb��A8�����k/�7�t�!��.]�P�}�9�X����{��w?�o���e%M��~��㟘u�ld)Ų6��<�5���p�u31f����S@�h>XE>�EfM'�}���.�l*|QϿ������SO=;m�����+W�����n;}|��e�o��>��jD�>�p��.,^�5���FL�|V��]s�z�L��F����v��D�������������ƛ8��#q��NT���0��11�CC)'�-Y��b�p;���l̽�6x�z����I)�)�c+Q�R0��˶������sPJ���e飑;�v�$G�Q_�)_aI#��y%��ƌ�hƾ�)�!a��9��\�d'KIa5�DGز�k�Cwo��.7�������MS�p:jMcp����L��&dT�92��H����t��MF|����\����S_�!�~ǝ}��W����^0b�Z,z�qJ��"����M����e�s���CZq�-�dA�U��cA���ͭh�5"�*>��V'{�W��h�P����6ea72hS��8gn!ƣ����c� J�8.D7u�v}y���`A֪��-H;�����,�|���S/�]�|K6���K]`�(v��B�p���D�bK_��)�t�8\|��H�Ȅ������V������z{�)̻k.
� >^��x�#���[���D�WE��`P��`�C���B��(�c.z��p�UW�������_����ǡ�'VhoO
��!�N!����_b֬Y�~�D�C�s�(�`r@�?�BW~u�%�9�z����-T�&��D��J��;�y�5�c�]p������|G���pn�z9N9�Dl��V�m����0���p�%�T!�5k��������|�M��v�T���)�����TM-^�!n�z���:�;��Eem/�]�K�e�E�/��{���[oBcSf]~�6�S�����^Ɉ����G����6��oӌڟ�3՘��,�c�~���܎$=78�!��3z���*f;�AMX��%MN �,p�7�5�@�=?n�!�*/"�h��w6�GCOьk��3��W���P*#��b�ݾ�SN�l�= �y�m<��o1hP���D8���/��
8�Hl����z)�y�o8�4
�<
ZeF>ɞ��̳j]457`�=���UϏ!c7F �B��E���s1�WF}&���
%�a���Ct�p�r�t40xfs���.hvNb4C��f���r�0z���73g"י�Іf�{a���(��q,���C��^��{��9��$f�W���7+��<��j<�G�Y��5Gx�����	XnKt���PX[�u-M�f�n|o�ԓT�5���|cq�Ģ����4���,�O�����x��J����&z:����-Z{ӈ�3���p��a���.S�C�2D|U��P���~)�C����FU7$Cp���}�N'�,�e�9F3|�y�z��"g,;;�P2��r�&��WKhilBKK3���/_�o��M�\֌d/kn�_�:D1�iX������#��C�Ǹ3qY�v���ڀ��s.v:�L�7:S)|4>��V�y�dt��
@Ut���J����S�_/�W]=ސ&,��B<}���	��A|��&�&{Q2Аm�.|h���z�.Y��n��ե������_ߋ�?;���EG{;��,�}��x��g��ɧ`��7���0R��Y�ҥ��G��WL9S�:��
�r�igP���m�>L�z�2I,|�,x�-\=�J�uwb���kq�ϧ`��G�;�q#R�>�{���e�]���J�ܖ[n��#G��g�!)�ɓO��;n���_����9���R���%�q�����nƐMGc���x��?��e�FX���P�˝���B�Ǉ��!'�@�C5W���xB��=C��t䏰��{�����W��A,�49�L_~񹒵���]ɬLQX	">��ip$�ʅ�"V2m.@$A��V%x�FC/m��!i���"b��̈|��	�S.ߤ%!�v2�\"P��c�j�ːDӂ�%$'���2BYZ[P��+��|H��WP����X��:
�Ţh�f�5� �a�f��w�@6Ӈ�߇�D�l�^�#F#�77�=߇=?��G��_߅T{14xq�pt����P�W1n��FC�U�Wh�bܼH^��������U�ֿ�UW�u=�j�k9���6vc%6DW<���I���ZS�e%����xE�YQ�(Eb�5&0j�=��d�=^_���3�w���k�hW�;�Ww`�#�EKw�4��X?���e���������W_�}Z��b��W '\(�4�����̓@W]�72j������!��1�0��"x��*|=�L;l�K#t/W���+B���P�*ۛԢ�ОY�l.e�A� ��yU��f�k��q�C(�!��H�D����]���Q*����q?Ǝ'�]!?��XJE��ɧ��������_�<�O>\�7�|�-Ķ[n��N��|(�E�>V�5k�l����ݝ�#hnl�Ǫ��� �� ��2���cX��b\u�h��)�������C�=(}丱�� ���/��Ӊ�:��J�� Ƭ0%*��e�j��($S�/��Ӑ�S��^��-&��+/��+���g��WcȐ�J�������⫯���Ï�T�Ͼ���zW=���9��mfo�K�|%Rܸ����S[����.]�TbDh��!!�ٍj:��������֬Ų5kА�Ǥ1㔸udR�7R�R�)Io>�Ď_M�8�ɜn�$�c!�H�+R�PA��-9�Y)#4��4�z{2�,$W� ��f������"\
�1x1��SFO.D4��`�����Rĵb�]�m�q�(9[��"�i-��uN�dZ:�"�1Mdʜe�7�MCJģ�o�T9%���)��@���ҕ�	�ѧ����1$݇A>��i%,9��d�h�c�ؑH��2��e9,>�����k��~�cԖ�b��Y�K�1,ր�/,8�t�P�E9��獕��~��tM���
~v(����!�X�6��~f_��[�1�6�`�=�)?�^��O��<�Oӭ,�!� YE���v8��	���Z���o݃�mi������=Զ�ՍۺU�6v� N�-9A�jv��\���W�d-#�Ǌ�(HsJ�%E3S��*�C���@S]=���2L.���.x�qtgR�"�#�yQZ�ꂛ2��r�~M/�b
/�g�W�N��@#=��2q��eik���;tA�\4����@O�\cm�����T�Ëb˓N���L�ھ.U�QT�~����Ïau{�,?{M�m�9��kO��N��rٲ�����_L9��o�&+���$T��r�k �l	�� +�,ž��ޘ_��h�"��ʥ+��?�G��W�vͱ8�<�h�� �
���f=W�v��Cs$��_|I�(�Iҩ��I,nV!/,ÍA���i�<CH�u!!f�ՠ�/���D�*��%ʰѰFt��}(�ۼ�*�eoϏ��fU�4���K
v�����Yd9,��W��0x��Q�2>_B0��W@	$�Ǆ���дa��&��$y'X����zx�Ԅ�23�	��2�I���]� LN@0D[�ZD"�F] ?���{1h��b��:�C�\�TZ�EE�3-7�!��xŬl*�L�}�tH�4� 헽M>'���`~�
�ndL6�E�!�&���$7�< ����:�"ԡ�p,��7�y�����nE1�B�.�B�����77�����,O������ս�w�=����m\�r/H� �H@EMԨ1*��5F^0"֧����Ɔ�ذ�D)i­��3s��]_��s�}��Q�>��{u��s����{����[k}����/�������,Am���a�Lo�[��    IDATN�G����)��ASGeZ銤5��]�����Mѵ�{~�5l!�����e�to�ҁ�J�����[��)V�¼�}�7Hq�Wy����
4?6��X����۵�]'_q���P1�����o9��ދ����x��_Ax����DN"=�F�d=3xO����PI�3gP<��)��X�����X��vBLP�����7L*�PYI�1�8�eN*�r&J���|p�WC�W]*-� ��l���w���KZX���>�$���V��eO�[��^��F�Xӕ��T,�e y@���4�c����/��^�Z�}��b!���M;�1����/���Y�J%�a<�D~` mZ��2��o��?W����.U�Ŏ�$EA�6�#���.L����#�MV�Q���&�~7YvMf34���9��d�%E�XŚ¥j�L�)!�=e��]"����%d�gקrϗz�#�Sِ�7*{,Z� ��ʦ]D*�Ѭ6�gG;��h��_ �}^ZdQ����U@˕:�� �L��1�Ř@(�3�d$���B Ъ� �1����Q'�"V��p�QY�E�����
�UG��`5(�Ȫ�TYE��B$���"� ͓�,�.{���ȥS<��+/��B���@VUU�kMe�h��G�`�4(��Fh��]Hތ-eƭ�G&�Rf��O��]�N��=g
&$M�E	R��R�q�R%�H�!��.�P���sP�i��e�"ЖE�d`����{n����X]�����:������F��2E��������r8]���'�H6&����F��xI�A4���=�j�m�U�����I���hU~��h���L�$�prɒ8T�#""���M`3����S��<�N����>���S��~�2qy�+'7<|��Z�@���%�{[���^fS�ʞc^*��$�@�c7o��w���.3=���(�1m��1f8C�h�$�X�����長=YH��3��ȧ�#hP&�uki�?���A��ْ<�L	z��l[�70Ϭ���-�}���#��&�@u��,:���`]��췼;_�j�4���ѬV�Wu��3mJ,��z�=c��k:&��iH2�o[����%mۻ鰴���iw s{ ��g��	Śt�U�o�=oFP(����ⳬ�+�o� @ ���is��z��P,ZM '�k�g�F7�P &�������$�b��`���*�؍6��B���z���IĞˬޜ$�]��iS���X����J��J��
UEz�>"Ɛ`�q��wĚ�Tf�r�T��^y�z����� �٬�n(����N�C�|������|~q���l�0<�c1���ȡYh���ο�
&����d�ɝۙ�u�o���Y眅v��G~��t�Hex\�i�:g�4�E%W�1��cP�Ay��h���X���=�L��듫��25�j��Ԟ�5I����
���4�f�-g���dP`6��4�Іb�Zc�6+�J�%�!T;-(�0�F��������"�����b� �X�x�<�yA3�=_���w��Y.q���-y��D0�<��-8�ռ���Ͻ�6�3|o���o���^��0W��Ƽ*�D`EGxd�� ׫8ܨ�r�?���#���rF�~�O�%�,|d�<��o0��&R&B�dP���E����t�lE�����d[������@E J!i97[������A��C7�B��`�R�D��V����L���D Fc8����..�_ϙ�(k�&�,�oԴo$1��:�Aq�6
���E�[Z�q��JXUu���|�k �j��B��%QYТz�`� ]X��J�=�*��P�F`G�u�-�~/�3H��b�x�-
L�&!���5����fD�L��Z��n54�lU�<"E�>d\!�hY��4ZMvcJE��K*��`J���CA���Z�Ȥ%"%�~4�%OUL"�f�2X����v��e��ӹ�J&� �A�]S�m�#�3��=1TEO�V*qy��L�wXW�"K:f�znF�X���[�C)��/����N$a0�M�=�dtZM�ʛ<~���)眃�o�����'aey=�&�Fp��`}}���6�r�8��s�%����p��)��s*��ɐbb|���6��� aWF<�8ӂ��K+�sh�@�L�5����!�U��*(���~�H�D���:ӳodm�R/��#��*�-�q��q�>�z�yY*��u=O[��¯
h�Kl*��2I��,U��6��MA[r!u�<m7���o ��3e�T�m�[Ǣp�6��Dϓ�+_��T����i��`K�x��xY)�gz�7-)���g^�k\��K�Û~ت����b�!�-�֢|���1Z((:��������p��2����~�e}��_#���rV��G7|FXZ|�>W�c��-�7s�B��hB_Dק�%Y|�Oe�^ɖOR�ޥ�eOZ��T�镉_������9�QH�L�Q"��;&�(��U��wtn�J�]O��{��@ �62&'���ID�27*���XdR�Jt�j�ˠ\�k{��ҵB���w�0<#lrF���	*A�zv^t��c/��L�mv�`]�IF��.g�6��:Ěf�o�v��rY��n�M��iq�jԡ��Q'Z$�Bp�i�����ǰ���i���d�2��AJ�]*%�� ���/R #p��1iRs�ot��"�E.� �8�4�=�|$]�Q�����\dI���(�A��!M�TZ'�6�;�H��V��>o2�����*/�h�� � � ;�L���K�޸I����M�K�--#��2Kx��	IS�N=�L���Z.����`͢+Đ�>+U,R;�
r'�������Y(`����|X��g�}��چť%��/"�� ?��^�#��
�d
�O�����F�BA�w�\T��]?�J��Ü�.9�k�|f�Y�{(��U�#A������Hz�T}�Y�SaK�6)CQ?��"�g����(h�._�9t��ػ�GDl�3V j>)�F_�9���~t:�5�g��M� V5K��ˤEAcҖ���F\S�9���")HZ�
d�ж�y��L�����į��/ɺ��T����5�$G�'B��}�z��ጹ�4D��M�=
½���=?cΔ{���t-�hܐb��	-}Ӣ.a�w0�B�6Q���_./~����e��G�_�@x�	q�7��uum��O	Dp���p����A�O"��A�ʠ�!cn���;[=�Jlc2�>� �⼬����0ɽ�$��ްt�C�ӣ��g�tä��Qu*��l¼q�D�#~=�}M�b��҃Lh?ۭ���g{e�C��e�wY��7���(���A���q�D2��jo��W�$ ����E�,�/�6�N��ϧJ@��ɫpZk�dN�s��-*��u]"^Q;���HjF:��
M�<SEM����J<�CuZ$�fD�,��]���r���8H2��H�c~i���t���9�4��e�ih~��Qo6091� ����:��r�,;3�������4��Hq���>�2h�����L���
W3�� ����7��T��������|~��Alh2� r�ǚ%�O��G�U1�����Ϣ��|����rj ��I,�/acm�l
�c�[X���,+N=�ܧ1����A:���?�67��cرc'��:f�����[Nm�H"	5���s$E�,�)Gj���6](UxdV�"���xcU��ǁF^z�"|e�Fi�ז�S����`eb�y��r���L�5��X�<DF�s��稂E-"�ϗ��� K�6�/Y	+��� �"(���=����P�Z�{-$�~��K��j�L�� ��Ó�=ZM��W��j��J�t���"g����(�jk��q#/��t	�gҪ�s�T�\skk8���pjx����>����}���[Ύ[�������;�c������Ј]l�������8��y�����	��Ѝ�I
T��<�s��AL��=�s���w��2]�^+m��7ç�i�.H"��E�5�n|���;[�#v&}Q鳷�����n��<�g5Hc5[-��bL�����#���&&p��}:L��L��"�E%�ރ+ .��� �ǫz L}l����bF-�X(K�׻#�T�q�i0q͆$:(��	ZGAP";n�&"����N��6�R/��iC&@��2��4�0m�>�g�Pi�Y��A��4�q$�K%�HEh�Z�U�|L�#�lM7�0� �E����l4���΀H�[�ݒ�'-�li�~�c��)ӥ� v3g,C�R��赔�6��E^�PfJ�Y�F�c �k(f�+]c��Q"ؑ�^ 27������������`�P@�TE"��`������P$�SO��~�߿�&����u Uh~z����0Z�O�>�`(�=|ݯ�X�g����p$�-M��Sl��e���
��86k-�K�$�� �H�}��7�c��q!-H�Ұd���l���.��|]̱uݵ:���ܐ(:MIrR��ȥ���ŕ��#�;-�~)�=�2%�� �,A��~?�7u�Lt�k[Ԅ��y�Ju� �wK���m;c�a�X���:���m��yD���$I�>AX����(�dY�-���8a6�j�$��DEf4l�C�M�q%tI꺢課L���́h*�i���N��lNX����;]���׍��+5C�]�/�'��[?�l툂�Ǝ��[;F�o�tC��K��K_��?Hs�'����o��O�}�?|ߞd�G����B�6��(ϱ��G�ᓲWr޺aӊ�@�s1�{�����j�r����T�Nz��-�7e,�N+j�L������~Μ{%7���Ho�Q	8.1z%p����i�6[[���x�B$b�`t�
���cA�*�ذMz�o/<�������:�\�ܝF���J��E�&��n��DA�|� �Jl\Q��ҍ��"��ҙH�m�5�-On���M�����$�&b� ��Q�X�p��d��V�J�2�f�L4�KS���@��2_�L<��q���%t-����3�,yAB:��t��!*M'#1��7Q#W&Mc�"E���9Vda�|	�	4�u$�I�K�q4@����4�'�s5eey�ߛL�8�_\�:��������(;��K�̢����}�61ɋ����� 2�X��q��4�9.AWu��ڱ�v�b���}���������{=ƇG0��"
��1�)~�p���p*=��?��P�]���L.7�Q1�+7˲KTQwt�~�Tm:�N?l	B+62p�?�_�˛�;�p�Z0���%�-H��AI�\c� 	����ܕe��(rC��YQ ��|�����_��>���sa������������v�mc"Ro"H����|E�'�ȶ̊zJ2�.�r�<V1׆{`遲yT�n�L!�#bS٘����4@=Hۅ�$
O}��xt\�q3~G	�q��#Ks�T*��K.*Cbt.mњ�G�i�R	����/��=�?\i6WQlɚڤ,#��-V�e��5]_ ��ӵEö�2eAQlEtlA*ɪ֚<y�����j�S�����Ӹ�*�H<�TK%)�jIm�_%+�����*�.�K�ӓ�e���AM��b��������tU�_U�IHą
��r�ReiK�?ȳ����Fc2���M�e�<���*�T��/��U&�P�H@H�ٕ�%�a�fT�*�b��x,��[Z���� ��2����2`���D"�TU�G��{�����T"��0����kgϭf�Y�t���y���^RfI�\�2����@ a_����<����116�c��5>ީ�	�Ӄ �2�������|��K��~�]?c����1�-9�����`.�=�X"
)���?�)��ɚ� ��,X�ւM�@RF����������;�z����-}����{�7{ˍ�����~���aw8mm����*�j���l�@�f�V��>��E�J�Le$�${=*�2'���� I���9u�~�aSK	x=fz���z7��-��ָ@o��7�C��-�]��`8��2:� ��麖e;�$��(Ɇ�ڮ�(�5٧��l���b:�{��??�;���w�o�[~�O1�~�@��va:�#Yd1�WZ�&����4���G����بV�ĮC$T��b�MZ��x��@w�N�7���ԭ#c ����`}f��Hm*�L`uy��2�N0`��y��������y�;?8 ��s/���I�������5^��xQ@�,T6��,� �T�N�R\B�s���x�睩�Lf�4G�ľ]XZ��0������ �ϭ,axp	=�~n4��\pj�:~q��|�?�)Oa�}�ދ�����8�N������옘B��D"Cj0��w':���u8��H �ۤ��{�&1�.	����<��K���'�w�N����8����ܛ�)�zh��ˏ<��	=4�7��SX�Ւ�n'hY�.8�$dF�2�u][�����!
%EUT�m7ֵ�ךLZ�WdK�܎�C�����"5J���RŔ�|H;K�$��rMt�2 �b��:������i� R]݆�	�u[�C4�/I�,;�NgI���󮺊�O���^�Ɠ�s�]YM	E�\L��ಒ�I�مc����E<GX0�������[3��2_R���U0X1L�d�'�I�,�ăA�W�5*El���OҠ�g�������R�E�F)+�T*����-S������;�G�F�`*9G�t�-�/0Si�@���i��J��;��п�=��i���ظ�����/=�YL����<����&�FX�уx���Ӈ���3`H"x�a���ٻ�+5w�y'b��6��p`��h5�H���d(�B&5�<7����6��w�I���$q$H�)�1���E_��kO����������?=R�``<7X�%��v��mG�(,��*���8��8�&�ڊ���h%���Uoq��J�M�t*��aY�ՕL]w������T�珂�c'���]F� &��N�ŜȒ�o�����W�[�r�[�::{��̵�XJ�XQ�֬�C�r�H=0���U��&ቨ?� J�!�|+�JfJS�+���kP�����ts��n���R�84����g��D
cc죺�.��S	�L,e�Tq���gN?"GQϝ�T��2�Nd&b�{���n�_C���1�[a�$=�m�S
 ���Yb��`,�%p٨6�K*�-!��p�:��m�A�����y���8����q�6Z��ln �����t6���裏2���e"!�H��P�P�ѡ�b���_U9��i~�ܰx����Q���x��w�s�����#p�F�����߭��|�U��}���)b���3�:�������Rf����Ag�"�F~�<���[i�f�}�Σ5R�"ml�T�4�.��yҐ4���H�#(���^m@�H&��Dkk<�J�m&����g���R�J%b��
� �~R��C`HYj�VA8�e��	�s� ���etʄ	�)3�Yg"X�V�ZF�Q���0K3��H�b�%xp��Y������0�����E��B��=�b@ߨ�����hu�	��&�qp�+_�#��C�g�dIYm�����"� ��p�mO,����P	���;��J8Z{�On�����-�#��.}����'�_������#����i@�m4�.,udf��憉J��0 �9͇Z]�_��/Hn�"KZ�.�n��AC,l��,h<.��4��.���_C*G����J�D"���)X�XB�V�@<�D8�@K%dQ������w�^+��@��NY9\�Vf���PVHs���t���옶��x�+��	�	�����pI�+�sH�#Ȥ��Y[es	Ø�����q����"�N"�J��G�������6����n�173�SW<[�    IDATO��s�K�T	uҪGx��z��x�Y�ԇ� �i�]�%�f�3cR��H��x4��c���E7�z���S������������%_޳��Y�p�4��ζHQu�	=��a�!����@�xW*%(d���G�4�E�Y$٧��3	���'�c�݆�m@�N5�M�6L.��EQ��Tʛ����$X������T`z-)��)��l��[tL�J&x	L�wʖ)+��.�o���^ʦI���P���3�o��afa�G��g�S���Ӈ�ǡG"X\^�)�ͯ� ���e��x>��Çcjl>I���<��).�g��dp�Q4�n҉&�e �SmduA8�
�&��مԛ�F8�Հ�|�������G?�������{N�|��Kޔ[ݼVm4�v:��dJC�`~�O��J(nnbll�A��͎*azi	~��ZG�D�]b�;h���Bb&;u�`��z�]��d���1	�	�Q.�xN�p��|H$"(�l��Q�]_I*	hQK��|��bs9���k�ʹ�T���2[z���0�+�.�-g�++�=�3OOOcdh�"cyqɛ`�Z������H�����<�Gỷ��3�4�f����0t�6l�-�e`(�D�kȇ�L�"���v��۠�ᡥ��j���#v��`�@IDcq��%T���F��mN�"Y�`�X{я�̝P'`g����J��G���7�>��Fڶ����lM5�{ր��D|�H.��:��$Oh��X��$�~�eMa��]4,��#�4�nut$lR�YS�R�VHu���D8�@�RF�VD8("�#
aua�gj��L@I༥`E�Oԫ���_���)�����>�zI�*�2�SI�2R"XQOwey����:tÃ��󼺸̀����Y�CO��`�p�ӟ
1�y��z	ۧv�[nf7�X(�}O9ӵ��u:|�����ý?�z���P��{��!��rX�D�woǣ��m/��Wbdl�����YD��	juH�T���դiOFG�QG����큾H���e�{}�}����z���>��{��l�Ŷv�뻩I8��g��Q����{�g��|*�luÉ��kP*��H�.,���t�مK�A�b�U`v �-��*���h(��"��Bl<r���M���d$�Y.�����Ҩe��;�m4��hO ��`LޭT�ެ��$Mlfc"[�-�x�V�8fffx�x3��Gc���X^X�)���q��?'��r,���A�/�%��Nq�|�#������J��C�{�17��x:��Ї��?ƾ�Q8��
�h�TbA84>��ً��w2cp*U��u�C��>�Jb���(C'�˂l;�EMEE5�.y�A��=����0}�=���.?��z�w�����Ǥ �]"�ܷՄJ��ޅ�?�B8�+��`,���ZD���uH�&t�0m#I\��W���{7�C��]w�y~|�yl��W\����pE�<�b�Q����&�sP����ܣ�,uK�y�,E�E���,e�D�"��̘��N޼������\�`4��do.wc�+E����#G�F����~.5����6 �#��?C�{5�,P�_��_�6�J �y�+�����W!�}�RQ|��������������r��8-;�T(��6���I�O��ɗ>�� n��]�Q�_�u'R����<r���uh"��mC4D�xº�o�}c�'~��q�D����W�ߑc�������h6��袆����Q�?�d<T\�K_�z��zP���-ec��b	�m4!֛,����������_�*\����Vo��mxǛ/ǳ�;>�9x�_��������u;~���cG@����Vc��̕��4�K�J�J Jĥ-��f��L���4�C:��0g�s�\�%w"�l��E�M�N����x{�h�Ã��>���?���u�ZZ.yj������;qΙO��>�wx�{ޅ��8�9��w��e<���ͯ=����ｨ?� ���bO6��'�R��v�_|�L�=r�o|��a��ގ�mb��7,�]>W@�$7�M��	��Cj��u��
�zV�X�/�m�#p,#��c������肋�M��y� X�SF2ZR �D���s�C"����c �DP�����O[[Ǹ�G�e@�� _U�B�Ɗ,�ɯNzџ���o�]w߅W�
��G?�s�~2�J����}��@h��ޏ�c�bX�QYY���H<�lf��R�M=�d"��UT��7L�"`]^^f�%y�����|���㱢��Q� �&�ʜ�\�N$9N��s(�յe�2�D☟[�$����B3����ԩ{��w��{�����=8�%/� \���s5����ܑCx��ތ�[���?cG:��_���4ʰ�M�p�E��2��c��!�0�"6Z�F��'��R�FL��촡h2\�AD�L�����w_.���s�\]�y����X��'d~��w<k���s���٫�E%W��k'v�����]w��QAm� ��")m��D8�������laD lXX.\Eæ�`�V�Y�r*^����������=oA8G0��G��>��66����W�-^��y�uؗ� "�˨��^ER��j�j���x�4���6/�J��#<7�H"��~�/,/yR��Ø���L��'���9O0 �"Q�󮒜�"q�yqn� #<2
�8�͗����5���>����>u-r'����K^�r��B�h6p�>���A4� �������m��N����N�U[��W��h8��g� %�pva��f��Btlv���!yϦ,��ٗ��q��?���'b��`E����?�<�WW�9����N���6L�F����A�;&���i?�4|�3_��n��3���.UYr����}��MDA��T�t�;�T�r��ȏ����׾�-�"����s~�~�Z��ꏣ���X_���g=��}?��W��ژ�d�'�ʍU�n�#�!���h5�iԡ(����Q���E����7
bia���*W�+���4L�/�������.u,���*!?±�f�  ��0#�>���9��*����`$����1FNE��� d�����v�t�0����&FG�p�zF��8���7��?�9lW�Զ	.s9xk�"Ƨ&q�]���_AJ=V���q�d�hYh�2������_��?���������������"��w����n�E��@��0	-IF���K/��{߄��|�?��FT�9ˊ��ػ{�G�p�u_�h 
��AD$�v	�|�{�ۀd�w1��p��߇��?�,o���n���>g�q��u��э����^G"�b7#bR��V:�@>�B�X@�Z�2r�Z�K������d*��K��[�����3�0�x)k&�**;�E_*��ꢷ�@��#�N����EV��!,�,#	#�L�Z���o4�0��H0�j���K���:{U@>����i�� ����� �H�^�`bb�R����J�趚���뫈�|�%m�]$�-Y�z��>�7%��~Y���#p�F��'�7���'����}�?�ᾜ�f�5E]AFݰ1y�S1����� ��2ґ8�V�e�\+��眃�d���Oa<�E�X�D>���E�ۧA�B0H5�AC(X/���napp�R�Nu��X<�`""	H�:�j6�E�d�Ґ�g�F����UL�N�X.�o�?�V�}H'�<�����*����<�x	���r�?O>��d���g��`qqR�J�qdv	�?�L6����Sq��8sΤ�X^]�����ή���#���b�&&��0���r�-U�%H�~V��F��@<������4	N��X�G#ҞǴ-�	��0t�����7fB/x��:�/�G�8�@x��/��+�.�]u�޹�w�U�b�a�2\Q�e(�&�� ����5�%�|m�C~.����z��h8�,`2`�YB�Ղ(�`�Md�I~����-���]oA�ƒ�Mۀ+;P�(����|��-��y]���@�TF�����ɣY+�y)�%�2�Q����	 	�i�7����iD����VD�A�!�49��Y֋p�t�+s�QO�0?�
�/�\&�E��l�޵��i�dsC�?sRTg���T`umD2l�
�
�0��V ��([&d݇N��T4�T$����m
X�(��0�s
Ӈe,�]��.��!��i(&��w�kR/y�g���#pF��'�����'���x�ޕ�~p��c�o�8@ǲ!�
�fN,��w(D�|>X���������{�R�G�T������\8&d���L��Vˁ K�ަՆ�`����iu��u��r���6�8餓�,�nP�8ŀI�A46txڛ�%�F�~%EfP%�&��t� y<� o�{	l��l��\�2q�/����G1��ѕ1><�#�#��AUE�K���~u�1�3a��47ꈆ�b8p� B� "���:��p�(q&�������	f�������(�,�m�}{�]Շ�����Xp�+^�K��UkO�,迣��#}�=>���^���-�x�ꭷ�4)��ڦ��с-:�B�i4ȱ�I��&��V�\�Y�$T���0l��� N�\H� �aA�}0m�&²�* ��>]C��r�(���D�� ��a�MOr�l�gy�� �����2o�܆"���m��YL�aa�T����o��������
###��(��C^�����Yf�\&���9.;����r	��b|h���j#;����Z��G1sd�H�t3�KȦr��ϭ,����bmy��D(��
�0<��(�h�6�ut�4��F>ׅ"
0M��m;�Ϗn.�}��l���-�S���~�Y��{�B�����G��j��nx4լBm���
�l�,�ir�*)
�6Ee�:���4�uĂa�Ri��Z�k���`�m8ee!�&`:6�ܶ��e@Su؎�N���?�V�	[�أ�ӵ!�B�������d�^���ju��c���(o�P�,z��yD�QDBQRʄilh�\�,��w�dMs����	o/KQr�h6��Ʊ���f���W6�"�� +ҹV��0�F�9�/�� ����3y�&��կF`()L2�%2O�IV�I�0�}-��z��.����Fr��#]a[I�ʂ( ����Lᔗ�|8q�e��W�я�	�>�_Z��x6���w�_W��*�v����f�_	��Ȱd�(��Xl�G,_��);k4����	MV`;&�{]����2 C���D��@���v��	`M�m@��БE�>� �m`$����
�&wlGq��f�#�U˨�Kqju���;�������2^Z ��2eؔ�r�l"�����<0����J����A���A�ǁ�ڢ���gU( ���&��Dz�e(-MA8����y��L�(,�@����,i@��!H:,I�����Ž��\��F�	?}�쇻���@ "UD	��UdH�M������q�}���'~��я���>��C/�q�/|A����n��eD�1��hD]�S5= Gձ�h����Lv��>��	����d�Zg�)MA$#Mǆ��X�#ȥQ�Ԇ�ɐ 0n�P$�"sF�����h�L�F�r�w�EauM��h2�f��r����I�k�Je��XXY���Ȧ��L*5S�K�-/�x��7�T.3���E�<04�j��Bi���X���j
l^p��:�|'?����i�	,�,b��a&�`bw.=���K�x�QtV����b�\@��B��J�It$eǄ�	����)���⶯}GD�0Y�$$p,����Bp�#�@��O�w�5����2���#p�"��c��������g�W�vL�#�����3����� �u!X$Yh:�9@L�Yԁ�������[�CVP��ܖ�E׬�� ڕ|���/�k��e�	Q�a�hh$E�\�"�(ؖ�ba�UF:�C�Z��f	;ƶ��@��� i =�2�ms����ES�K�*/e�[�;�`�5:���\��ިad ���3
:|CC8�qɕ�s�,/��o�)�H�ލk��VLN���^s�L��0�@E�{�Ʒ?�OSDL�2�YY�f����8�PKfkFO{�E;i�t:� ��o@sv�f88.$�#��ħ�8�df8�̹�8��~������O?�k����F���>7_p�C���S���w����UT]u������8�I
��g:.���$e��*��
��â��cc�S���/�c ��������]/~.`���Y\���Cca���U�|n��ǘ��t/��w��8���ӿ 	��<7��bpt�z���;ƧЪֱY, ?���*)T���r�n��֨syyk���w�|�lG��x;�&''Qk4xi��	T�K��lBF�ԝ8��d�����/a$��K��|�3��
��o{+���~� >�����7��L�[q���D,�=�Z�U��5���i{��x�����4�8������������ms^ _^�Y�M"�䧞u҇>t�	B��6}�������ܽ������HH
Z�.�`�BյQlT�]����?�/�{����_�a��Z)QF�kA6,﯉.|'M�+���F��¹{΂���5�������y8r�=��羈����~�#x�;��u���x��O�o3P.�S/�3i�Eem�5�����颰��]��Ѭ�Q�XGv(��b&[�'�U*h�Z\R�r2�,��4�0e��r���ccc��6j5l�چV������(oj"�Z~ ���h�@W�v��G�;^���a�TB[�pֳ�������~	�~�`ߋ��O���1鸘Jİ��K��u��������_��(b����(H
FCI�h�8�U��v�{#Z2\h�JKAۻ�٧���������S�����m�����7�����^�m9��W	�٬!0���9g�(��'F������߁�'������Mȭ��.NNd�)n"`�좕M⼿�G���? K����W�n��O�cصs
/}ۛ�W��x���Y��s���/5�nO��|<�Ig⃗]�ݩ8v����P,�al�8��76�8e�n4k��� 7���f�k!ˢY��R��Pe��Կ%V31��	x)�eQ�j���;�S��Z���P�J��r��q�Z�>��0]�'>�!���obci���Հ��[��?��j���wq�3/��矃O��2�R$��#X__E��A� ��|�ؿ��#@��M1_ Cz������?GX�aT�i$�����D�:��>��_zS�t�G�D�@xO�o���O(���\��.��R�4��lEF�4������g�'<�������;PX\CPձ{�4������7�m���6Жdl�ڑ8v>�B��̋`h�P]\ć��{v��k��+|�����{�� ����O~
�w����⚗��$b��QXA�YBf Ϟ���&��<�zK��񮖊pz�۪�Q�T��L�-b0����4NT�T�lE�e*9�L��m��+H���t��m���h��x�߈ǪTMg?����b��G�k>L��7�g��/��(x��;�_�����v�4�%�(��X.�P� 1���핸��[1=?����~�A$�L�Xy�!D\F��t0 ���H�YQ!�+<��R8��Ϲ��/zB'@���G��q�e�w��E���o�����l��D@.�R��A�v���ݻp�ŗ�?�9��J�&	h��n� u�;.GR SR��b�Nl�#�M��,���A�����׸�O_���z�u�x��㱄���    IDAT�݈�t��Q\}��kr/�����U��rl��P^Y���8�e���ݷ{�&f�g�%9������,���,,��ɼ`px����w||�j�����8+&&� "��+�������6�#�8Rk��?��1��������_��=g?	C���'>�O
*.��r��,/��$����$"a����e�P4��,#<�G~jS�����5�{�]�U�p660�h�ڲ�yjˆ��i7�5��W������cw���܏���@x�m|�[?N"P�����?z�҈��|�.l���Iп���*z6��� z� B>?:�6{����mv��F�Ttj(���߶���E[0ZH=�8���*� :<��}�K8��`}fl{csfmel۶�tl۶muұm۶m�c;wlc�y����O8��^��1��-�������3���l�j������7F����:�a�������V�ֺ,�`��3^[�T��]y�9Z�~1���ZS��Hɠ@-��=-Qf�o�x�gzY;gO��1q�oR;��##[��~�R�i�jDbI�*j��,��C-{��O�~�ҩJ��Ǚ;v���މ����Ppȁ:s��Ӝ�pT8����7v�ؑ2X*f�篟,�+!i�f�z��FV�<�(������];9[?y���x������]G��@����W�1��<{l��,��<�߽|��=���z0b�Hk�~z�G6���k�8	E�f=��_Шe7��4^�Jt5����1=�i�q���Xء\�����8A"A��j�j�1���vF4�>.I���l<�#ޓ>��1!�sF�� -��`��m�4	U����`��J.��f�t޲�e�vj�G/�F���Z�I8�%Z6�
��b쫦�v#���a�Tiȏ� .�j�&̘�:/߾BMl/�&=����m��X�ӎ	���5�wQ�B�+9�7Q"+̈́�pd{I��c�:�c�C�a�D��Q�n w}f#<	�_:��k�>NE��<�zn�	Z��n\��YX:��1O��i�>��z
��2(��T�b$�օ1��3i���|�Ci
���4!�������K�hVq��sl��K�(xZ�@&HxH��q��(`0a��1��g�ţU�U�M�*Q{<���T�G�p�1�<�Ħ3k}\�w�����dէ���+��emjJ/dq+������Ud�Z�7u��T���Õ���3����E��O�v������5'I4i�L���B1�6H�d�srr�%f7k*�aWR� [�o��s�H�z.rlܾ����\�����v��t:xF�a��T�|j@>e!�?�~Ϗ֛Z��gH"�.�i[*AT'���^�))�
LM&;��8J�K+"���5"tmn3�������ؓT�y�A�7�FH1�v���3q�3�lP_rG��Z�Ag0�&N��P���4g�GC���]�1�L*4��d���Op͒��d�ܚ*i F9%�+id����ƲS��`6�J����Rza���%>f��CU]K���;Ԧ@��4o�h��6|�l����cE���n����34p�����,x��lǒ�;�P�r`UZtU7�h�;�*Ep6
��2��+M
Q��x0sۮZ !�9k�}I�FQ��� �^�������p<ͧ��'Xq �˦��.��������aQ�)�`A��k��D�U�	�-6������_���ʲ ���c�_��qh�h��q��E�{�-�^��T�����:�dĢ-Q~��u��-s����I	�Xب�������`΃��nV$*�֩)*1�hΪ��FUٜg�����'E��8YIK���ߓ3'���I����u���3��G�x|��+��jn���	�����GBNs�؋\?�"1r렓;b�\L1Co=n-&{����%�w#��)��,uqԃ���?��ձ�/@��9��-��P��������ȄP���me(K,�nQ+ը�Cv]�h/���x��������՚n^�Qwҟ�=v��l��βp�d#�wl�0?_���X#�g���gb�GpS]��oك��fɧ�Ź#6�hqx�����]��*<]�ﰦ�\�
)G1I��{ǖ��z�M�����n����@�/������e�F�Eϩ�ˬ�/�q9�XU��Vs��<62S�.�i�.U�>]f��L�mq����YF��5Yb�ig��O�o��� �`���M@k"�㞈�7����X�7.�s���.���'��!b�o���舙#09o���9-�(& ��Y�U�G�b�m�vM���PY#$Y�z�`��!��x��J	/�N"��zw�M�!��t��XP��%�jgo���j�tS$�+�W�t�mW��N�ڴ�%����p1n��7yދ�@H�_�����%�2$�`��2���M����DZ�2�UR����Cc1�yW0S���­P^ib����@��Gnq���a��Aܕ<�_q��`.�N�@�T=<(c4T5�R:fhk'�twv�w�4ٱed�a��3�q�B�������ki�c0B<�э���k4H �݃O���5�o�y;�5����l�?xNSѻS�]7�dS�ZLt4�����gꑼك���?�9��g�䱱�bY��ؠ�hj]��ia?g��6ܶZ�\�K��Di�M�C��{/�$������d/~�u9a� ���Ү�����o�u"+�X�os�7/�m+�[�Ѩ��Zm��o��������b�s�Q�:�]3�%A�Dq��1�M�q/�r��U�P*{�H��u̧��KzrΆ"�	Ĕ"2�7����7�{j����[c��h�����m��"��b�3BB�C%ھ��i��lu�Z�x��[A<�&�Y�%���O{��m7�AON1 �Ph)Ǌ�7oy��o�o_��v���X�h�D��z��}�4JD��Icj�st5����}!6i�8Cن>E�m(f�M-����T'�N�(���������|�ȳ�,Ϟ����8~�U��Ld$dK`|>b�'�����mX��1����*��H����O���!�_���|}�f��/��+'�?Mf�">��`��W�P ���S�'���QH�%���,6f߻X$&�VF#Cwݎ��e��O�4Er\���?UW�wBR��*i��|�X;93�����(�`�R"\4�VPo�.�� cG�P�E� /9�Q���OÓI�9��+hv�8PV���^��p=���Z���(/1�t��it�׻R,�f�������(�>D���K�Oʇ�.]���$d: b�;&7���@9d&|���'>�nh��T���#ό-�L�z�&#�%mI�y Á�V�A�HK��%��i��1��aڿ���7�ڟ����1�}8��Ք�U��n7��@N�1�S�`�.ɪM��r�S�T��?�p.!G���`��e6�����VTA���Y��U/�@��_���oW�#-Rm�!����-��zo�y��	��Nڗ��ޫ���ʔr
��R�hml Ka�x�	2￉�
�g���S�E	�����rI��	w��9����6r�Mh��"A�c�s��}��`B]�]"����v��w�ꔟ0�������w��߃?��}��ݔ�m��wFf�?K������̙�T�L�oJMuCb�n��6+M�Q޶NH�m�6�� ��5��Q����.uB,�K��DO�i������BC`sA���O�tdg�<�F��d.����g�i^��h��e^D�VZ,�z�:2u�w�y K_�ƈ�(�,�'��R����E�:5������ڸ���q��An��
�85Oo�u�|��++�U��0 +��=�f�Q��_?�i�W���E����M�B>z�r���'�6�l_����O�y)6v��v���SU$�pw��LNN�?��xX���;�f!}��	r�����-T�u��t'/�9�\�K�}
����$EOW�A�C��|R,�܉��+_��� ������'!5��Gm����9�
\i�_�,s�yׁ9s��ӤkBs/������M1��X��V�85�D��
�m�Z��N���,�@����7�y_�?� �~�J`��T�X52obDp"ǑEqڳ蜛���0Y�"�d�R̛�����9調o�#U+�MZ�����>L�b U��7@�"[��������n��F�솤�ւ���jwh^�����U��_Ԉ�f�ǆ��&�����@�K{���?���x�*�Q��?�g��$�2��T�Fc����3{@F~��@�4ߕrL`�Ō/T���s�2 ��m�vr�@�w+�,��Q��������x��N	���/�����d �5f�>0IW_@<������+�8�)�����Q"ƍ�����%o���3	�<�M�fOO����;E�ǉ��!�'E���m�S������Y��\JV�Aze��*�lwF�ڮ��eޗ����OP��t��	4�/�e*G6`���j�9����RJi<!���?�ԉ4��d�����i�)��i��[")�[xv���;;��A���{JNz[��	e�-�}�c��(�<�;ڳ���g��wٹ��}Z�c��S_/Mgo�Nsq� �&9�A�؁� ���D�k*#+��/�vj{�:M����t�7B�㯼���p�J���錠D���%U		�qg��?HH닮��#��~���!�&��Xy�'���K�ts�
��\1x��z8B�<w�ۇu�&��P�)G����k�tß�#��~���5�E�UX��s��P�}niawB�i��W-�<����=7���Zݹ��B��"Aba�ZO��
���K z�J��묒�%�c6>�N4���J����U�	���3�3:����5&�����y/w� ��SOW1�����4�<eyjT���(�����cܛ��\���<��Zf�X� ܾO�ڟ�:&ל�^��پ��4�Irq�\Q� ����V��%���9�ISI�f\�{��w����Z���r"���\�o0���O�Q���q+�~t��p��^��!2%%�%
�M�[�Ya��*�T��sGs�+	1�4�h�ϵ�A�I�Y�[���i�jF6D1����~�}�U��:"�JL���CMN-�j��3EB�:���b���*�����:���za�QzTrU��H����Z�ʀ��p��$�����[�١|�$��~���)+��4Z�>��P�G\��<���0N������I2����G�E�AW��6���������ί��=5�۲h��l��o���x��㉜���f�n:qLn�f�x=?�(�ݫy��sEE�*E��nM�!��q�l����:�zJ��7إU�S�Cx7ЩՌ{��ގ:�yQ$	�N���y��\i�J����R�"��im|����vL�.�I�x ���s���c���]��<&�\���G[ƪ�R10���p��x�éy��-'�d�̗�C|���-.l�̬�
f%�7v�����T��%T~"�i(Q��PjJ��ͽm�)�lv��i��߯޹5]o�$�s��gU�<r�cO>�%*w~瑣kJc{:J�}�����9Y���`y�lA4���Ow�T=�L΃N����Ǳ>oW-}�r�k&g�X�q�O=*xNG<m�N���NKn��'�����}}9�~1�,A�K�tt�3Ŗ
e��۩I��_�X��IMCK �byb��@�������`R��* _y�F����^�P/�F����e�f,d&V跛�èR�.��<�dX��
Nkg\��.��kwI�d�|D��U�^u�bd��mRu�\)Z	9��T�R;Z�
X4&�V��=�|0�Dt�-[0<ڪ=0�L��NS�T=�m�]l�Y���+J��M��:�A<�`rJbf�o`��@����Z��2{#�t�'�j��V�W'E�&h!j���,5��f�Uc˜ۂ���(iD���t����ݖ��T�r�a��-r���sr�SKK�]���$4s3Hs��f,2rs
��$�9���R���$��]��+��W�����F�n�ͺ����ml|��:y"�Md	��s�2��rI7ץT�5���dD��	��[cb��a� X8�h��S�Ĭ|gJ��%k{rd}b+B��C*o_B�is�W��d@��?Q]&��e�K_2�c(I.�e��C��,C�e�*	Mӗ]^ �è��~��϶b{	�h�Z��'��^�ĕ6Vs?7���M����kd���P�鉷�rMbxQ�"��o�ݕ�^Ei1W�c����L����8��t8�Y�T��� �\g^�!�A�}��umMҵ5%r�bz6	N��ŤL�(GBȨ��ܴ8��"Q�4�?��@I�1dӖHF�>p�1�+�-v��E��{�l��?�0]�^�UEzJ�(��Єi��3��8�ZbI�_?rT��s���6�+"��`.�4*��Vr�0�v;�>�ʂT%�׏7	�&�b����"��L
�Ռ$�����N(Y�[��1{��>�I
�\5��L�[�:�7�1%�,���)щg���G��sw`�#\Iv��g{g��&� �Ĳ"	EA���Jx~�Fn���xn%2�0�Ҹ T3�Vs��}|�]y9�y>j<���Z�g��l�Dț,/7���$M�n�&���7�q�����U�.�����	��z A����3Vt�z@���Q������>��.H�@Ek?u:�v�}��+tçx�ӏU�����qq=�#�)�?��[��Yi2���Ue�n9N�d`��}��LE���7
=�P����ք�,3Q��1�F� �WoL��u3mc�{)f�I���R��0���>Wz���R��2Gի��k婅��@,����.8��&M���S۽E�Z8{'�-'QM6j��.�7�R�� ���H��2E��4� �)1)�M�1��L��!�,s��[V$[�����l	9JJk����S�rQb���r�V�|k�\���13K�������
k�㓇	�@̛X�W�r��ȏX�k�d�l)Y���z ���ZxZs��_Jh�*�aj�%��t�gw'C/�gۢ���u\�B$F���2O��zagY����H�[ߴ|����Ji3�9%��J~Oʢ4����л֕�Oμ|�!�H��6u�av���u�J1�SM�:���4�Nhax-5�Vɋ�yO"\��X�d�QL "b�T[J$���C���
5�����(Gf����^�Tn7�Ze��H�(��)�M�dM܋�w�P�a��T�<+��4�Av{�H�|�9f�d�L���4]���'�$���EUM�9<N�:�0�@�k�����@������)���S�$K��LAӗbr����G�����5��t�'�̯LS�>���6�"�<�4Z��"��q!O��b��p���%�OD=>V;X�Ҟ�l����<ڈl�S�ۤ�U�;b�/����hJTc�A��R掺�@X~���q�p�|�h���i#{��%ޡ�g�E�V�&4������i����/"l��n�8ȱ��4���ٺ)*+L`�x�Bo����#IB8D�T��m,a�ׅ�u���x��M�CE�3�k"E�Dg���4m/Kƶpv��O"ʑSJ��Bl}q���ފ�O�i�j�����a"W|Ap��, ��˃��,�%WS�K� /����~s��.�.���!�_���Q��X�j��htǤT���aeئV����fq�҂Ct�+~
���o�T�W)o��L�V�43#im��F�&m9����҄W���>�U�]L�.`��cC���H���ШF�@6�Xs̏���q��x^��rW���_Q%��{���V�����>���Y�_�+!�qx�Bq�k�l���@z�fMک��#�Q���N���E$�:E���D<�W��2�Wֲ��C,b9���P�d��2�}���Kk�g/�����u���,�!��	����sR{��f�VJ�>o���MQ�f΢��l�
��Ӊ~J�Z��蛅�t�Sƻ"��'���,���Ua��H�k
ᒲQDf��j:���{@�����EA�히6pvq1����D�i��ŏ�wh�i,&W�~ק�g�XTCS�n��	4�(��B�A�a�{>��Y)�T�/B����8bB�K�,Q�ꆩ����y�]=zp����F����*qcm���/v��3����
�P����+jk9�  ��lw�N$�,V�d��{V4j]B%�(��=HMV�оZ ��88�7��al L|�r�[�0�%Ƹ0)�*0�P�>�Aƥn���o!��ܦdU�P PvX1܋�B
�M2�,�7h�:D9�ILt�3�W��O��� �!d�@G"�f	w���I�Th��>P��\��ۗy9䒥X�_h��ď/C;Z���e�~�e�W��<�t+e�f���r�Ɛ����|�ӔqΧ�����n���OzT�FT�+}#�S�Q�����)ߪ<��U�8�	��5�n|��BT��&����ՑG�$#$UG�Q�=�a��=�<u8��#��TqMn�?*`���Eu8�)y������ǒ���N��RJ�D)�%���1^K��H<#U�1<J"%G���H��h�����P˳w ���]� ��{��Ԕ���P�u�������ٽ�I� �!�ڃ\��O��XZ���>�[&�4����oO��;��žA˲����T��z�����Eҽ �h%��`Ŏ{����$ Y$�G����e0?=�n�������^������1H3�}X������;��s�l���c�Za,9Ŷnm����|�%��eSjߛ��������-�*S�Tl���D�#I�^�IE#&nq<��p�z��i'�+սb�P(��
�������7�l��D�0�o�lQ�����Vhx����Or��-�囯��k�y�Z�����%0�	���QFZ�F'�2�?��оTbya�s�ب(6^��ó-q}���7�h�da���>]>�X۝��獲�'-{����M�}��AG����7D����'���|%��v���5H�`�1����e�����ԭJ�*��ݝ��I�Ft�\���d�b�Y3�Ȅ��� #�u@;��xS!��|�S��{bi�6?nߎ�~���r�o@%�f���X�mR��o�G��"���S��R9�}s�����
���B��if7 ���4[� � m�
�`��`DV݆N��-���sô"��E�`,����%�k2�Uq��$�Ș�%R�|N�*8��{FD�&�>�O_���n����<��u��������W|�,RY�0}(�4��'�œ��N�u��J.�i�*���P8��n�\O�Ic��������|��2����G^��g�������+�0}��������]�I0��@�% J����Q�:�ڏYt��)��].�d�	��54�J1�#IJu�.�W�?#8��ٳ����C'�!9Dg�9x��%PO�{�l���`��,��zsp<��h�b�?	���펑�>��5_�6�����z�ڽoL�Kğ��%�y��㓳�3��^t�0N^�|�=����f�D4�F%����95��F�)���JM r&Ȇ:�>��R�*��r���� Y�b��7�@�����z��aOͳ#��@����F݊%��z=/4VmNOt5@��*��\zo�/}~k���_�ܩ<7T��Cb&@�/���+ꪑl��3v��W�}ϧ~���_8�=x:m�b�45u׏&/�\��,%x	�q+�rL�=~��|����0�ޫ�ˈ�g��f�t*7.�t�Chjg�&؋)e7?a�F�W��6Ǝ�՝��8���/���^��觕��A��Wr���6�k	?��������Ft�:��4πx�7�	�n8��͙ �inka���{{d�������<�cVO-�����|�����2�i�Q�XWe�9��ֿ���s�����K��Ts�A���_�a�u��H<��xe�ɴ`S6qQ5��,��O�8���O݋�����˄�������r?�}���������5(�/'����?���+&�d���m~Nҁ2Vs�bg�'BѬHi�������f�$�P,������aZ4��^Y�Px��Y%��]oL�2�������3H8���3���|��U}����9^p��+�f���9ņ��ˋ�ؠ��Dk�k')t<sp��J��d�cם�D��K�@?>�e`Ԙf��$U�~�K�͕_Xf���]S�؋>���������8�-q�M1e�������p�CX�y�|���x�l�\����� ��sp������\{x0�r^Xv�
�J�E�9���;�0F85Ӷ3<���y��$�S�D�Vlΐ<,�Ph�M�WF����~�w�K���o����w��*�5�q����:4`W��Tr�}h��iaak����I�z�,�Օ2�`�w	��#	���[�R�E���*��{�q��|����³4`U:�Z���B
��,�s�>��f��|���ZY*P��z�ӿ��a����>�-���KfG���F��㌈6�A����1>%��
).���o�S�nf�>%��Ǉ0{���z��X�Jzώ�E�1�R	���Z?[B�L�bɶ�~\K�h���[���g�
��� Z���Tي�����P���uWu����K��+D2,wi���Si�P�����L�
-��Aq���u����R9\T�?FzO��ū��c�CU������*6z"��9�[}14s�+�齱���p�l�gLL,��T�[�����03G��E$M�Ϫ��M�p1���Pe$bF#J�܇^��y��dJ��-�̥�iX��/�y����R�����w�Ig�Q^n&)��%Tl�'��E�"t���lX88F^v�#�HR���x��
���.�8!�{��?p�WW��uu2EABo9�=�k�DU2Q`���%r��mv&�ޡ��I��O'4�o��3��XL�2nf��/)�3��=�S�Qy,��Pyˮ5�$W��'��ʘ��a�Bra�%�b���*u	�%dI���05��U�AlpSc [��r�� P�����-hQ�gm�똡~� {�|ߤ$~̷�8q��&E
t���P߄;�(R�%��k�W��o���Z�Sb=S��Q8�e� �8UO��:	�P3gsA;eT�������[:���z��R����J��L��y�2t��L5 W��6*!+CKEiZ��0	-d�rd�Ti�>.F4z� yR�_���zt�L��G[�����!��h������������t2�q�w0�Ι�V1�Q��z|ytvtC�a;��c�W{�����d�3�pG��Cb5�
�"�2�`8"U1kR���x��'e�n�HPKX���4,�qo��M.�ϩ�T/%�Be������*r���wJ�{���_��Br[�_���`�P"$�����MIiH�9|#T,W�5�����$�Lf�:���Q��WWlbOMO�u ��p�<7���9�� �v��Pwd�ȖMJ"�Ș����f7���,U�"���.��lqyg��>�
��ĬB�D5���<�`�Ԥ��V�\9�-DK6��]ZKJ���j{�s���=V�=�h_�f`|<̢M�·؀�K�jq�sX�*���OÝQ�������f���8٤�.��+��X�VfF�o�������|�*Qhjʊ`s����i���ܦ
hh9p�a��u�����3��?�;����I4�m"U8����.������{���nu���	���ۚ��@1�e�Lc�6��%�	'$���\Sv�Ljۨ�Q�W�"x��H���bQ)%0�|g�+o
��&Ř��SVH��8���xI�������g���׀U.��d��pnY�wp��%��2�O����2
��܇#�����b�B�������o�>!��8b��%��_][�P��TǮ��c�_���,f��`55%��B���n��X��}~1R��Fe�xikѴ�O���I.3�<��	!^��_�Z4V�Ic,���>u��B��6Γ��Z=�	�`?��җ`�2wI~����u�w3��>�ٹ0��ߦ�{g�d����X�6df��Z�a��k�|�h��۴T���#�g�N]�������M�c����YTk[��Q�b;�|��Xc`栘�H�ޒ�j��m�`C(�'�͉����9���c�W���MȦ�k���H&fH�����C�$��_ϑ'j)�VX|��	�`Z��n:��o�[1�M�y�E�CEF�%��L���=Iv����H�s5��Ss�1Y�N�
[4�T�8�f�eӈ50Y5b����� �8�8��pa��x��L{�Z���Gf�yP�2UJk��f�\�=�tj�y�)%�˯-�ޯ��o\r�ՕSP8Y����[��K����Nꯒ0��d��, ���q��di=�%��6o	5�X�Q�m[�=�u�m����98/ #)��9�x��b�^?1No���%��L����µ����r��G�ڱm�N�Y?��3�R�N�c5��acc�9�k ���PĈ���(?��ֻҠ��"H��<U*8�2=�.����m�x�҈X5U�/�+&�����j�����l�7�.��gq�Pa�η �vh�"�N�uh3�qȠ����_ކ�̗��80$�W�ʁnZ!Eb���S��Ƙ3(x��D1�>{���c۔����7Hd��%>d�!ŷզY�֙�2��x�y>��L9ܙ�}Z�ʔ|�(�o��-v=�G|d���Ҫd3W����R����9�!^�j�U����|�e��D8WW����1Ս�j{�4c�ژ�'5�.yH�(|,,S;����Q:`��йw�ʩ���Q,Wgg�x��_�kQbR����)@�࿣�7Zpe����WeS,{u��ԍ��JA�&�n�R�cBF�yxx����kۻ�`�T�u׉ƌf�� �"�9�������C-�z���gږ�Ũ���ىC�	"���Q�|l�%5J��ɍc���tJN��xn"o>�����-����wybu�γQ����y���c:�a�B����/�)@.!�tE���L�l�'b^*n���r�h��D9�&v�b�y"�]���b>o�Sԩl5Q�9PZ)��h��ش	��B�rM��U��|�xMS�T�zqwshc�&F;&��(c`��LR��N  ��.5?7-J����ʗ�'�b�u��)<G�[F9782�����/P5��?M��F�����c~]f������j��d�����b�Z�������:7Y�;agb�jA��};>�9I�f����}qM
�,��H�sb��5͒�n�*��|���-a�%4
�q�vh��f2=�9�����[����u��y�1�����]���F�#���/ŧ����a4�Q2��b	"�/(�f�3d����=^���<�k���s��6TC�K�V��&����d9q�6��M���Y�6I��C��H{>�C'�x0�)�<�G7z���00��O��ä���CB����f���N��.���J5�e�U���^���XE�i�G7[�td�0�����u��1�0�-����W^cs.�N�1����@/7:�8;�$���rt�ŵ����|�vf��;��k,0�^�Q:m����ow��|���m�(�L���@��*�Ќ6��͑g�U[ұ[�����]ю�7�S�ä�א�Ź�u
�1���D�>C�pC���l�>��ʾ�{P������C���ڷ��4²�J� 4��d�y�g�Thlڜ�J��XL!��}�6�	�ኋ�5L�)`}߾�6��'�s���w�kfuۑ߂����	��b!�0(��*	���߀:��������%��o���AQ� �Z�7x}lttCgk�]��˓2C�m+M���x�bB?m�A����o��=��*�`����=��^HD�b͊E��?bsFM�c��F��/��YǗ}�<���y�l7^�f�=_[�S.SO}��s�i=��h���)FĻ@���:����W��\>F��Z�)�f�L(U6�HEJ���kֹ|ӳ�D�|��Y���w�T#$BF9��A�5������ � x�OȎʶ�͹�}�-��'�-3�,�|�|J��wU����k}W����E纒�	�v�w O�� h�`��q9"J���ᅌK����9�z~��n�g�Wz�������ܟ3.���t}���q���]�8����Qc���hj��p��g��x5�4M��r�M���MLPY��mn:Z�K��.��d&S	A�*(�}֎G{\�O��k�f��i\2�w�D�ak�W�Zy��?����A	�ߵ0J��`�~}Z���A��������p�z����:Rcl��{�wEx~X����j�2<x���9��>�q8�L�v��	/�s��eY�SC���;$k*�,�y�)'��N%<���-�M��"+bY�!)j�-�Q�;�|	x���5,
[^���'��������AV��Gn�z�P3Jc�S���֠�p��f����0b	p�+8� �}3����9�51�{E+�Iԥ4챼/؏>pi~Id�vXv��y�ds�{|V��Kߙ��o3[�3-� �_�w�p�Ϸψ�q�=�o��ui��<1�w���ik�:i�uT���,\|d�4q+�f���3Ԇ�Qr�Kw��o��%�qMZܵ��ɘ8�x4�!��dV+"�{��;wӾ=���i���m�C�&��5�F9��cׅ׻J�d������C�ٟ�����"�0ϕ�ܩ���s�����hJ��lK�1������+�k���=�P���I,��MԝEN'7�2�J����H�h��ֽۣW��?�q���
�5P� �{!�G�#�,�ש�wt�M����H��TϟVi�-�>drT\&hAɹ��؋���-��7�{j���u[e��lc��RL��E��72<A�taƸ_�����{'��=�����u�>�ݶ3��j>^��2eg����,���ysLxr"�hv�����FVi�d��ez�{{�'S"U�p���R*ɽ���n9�ݴ�1�iY��i��+E�4}B�S�L����Oi��^.pq����^���,��Ut_�S?��c��L�-6x�r��7.����pm��f��:t$��S�f�>��U��Qۢ�����2�����ǚ!�?T36��K?�v{��?n�~�q�9I]fĉ+{ݑ��=��#�� zPXb�2i��d�Xb�N9���3[�;��P���B�gGM)V�?"�p��4���Pj/5��oc��hn����9c��Y�k�T��n�4/���/��$.D��8f(̱��)u������@���l��M�G��������F�[t�_�COJA.A��1#�[�	���@�N����l���$��P��~� 7C�V��Tb!X�u��i}��,4.vʗ!p7(�K�X��Uas�Z���K��o� 7����͵�-��q�Ӿx�����Φ)���]�]#?�?-�<����r<� z/������c���e��w`�Ϡ13cһ2���t�ô� �[��q�L��t^��q�Z�6������8�e$E߇Q1«��U4�*��&�������vVb~�����C�������J����ô��ȿ0ĕ���ũ�I8�e.cF[�ۉ�l<L�/��h%�W����H�Z�?Rm��Z>,�|ǋ߶&��#�g����T��w��Z�?�����O�On:a=��c��\(a]X�F�!�6�ab���nzؙ�Y������SУ��'���dԄ<>�I�%��G]��Z��k\����f;��K�ѥN��ɍOLTqi�CxQ�FSO ���k�ʻ�C��'��6)o�2:�åF��͑Y��3���I��#��B����w�S��'ۨ�diT%D��'����2'!��?��m��yF�%uv�d�u�0�)�T:��5`�G�+��ބ�`�^�2�e;N����n��mh��;�Ȣ�Ӷ�(7��v}��{fYb&���#�.k>ETXY� �<�t�"^d�	L>��/3�w^W��pF\����9TE�Y5xp���%y
ٮ��3�r��XZz�U�vsR�\R^�&MKO/�_ظ��VV6Z�$ظ�,c��B����V��-ʩ�4�O�| H�\�)�3�� ������DδY�زs(�ӥ�D������~�;.���S>���e??=.���'t�rd��>6!G�
�*�d1z�]RE�jK���[�}d9���3Ȭ��k���xQ!V4Q.DV��ro���9���?��������Fz��?����"���P�Ќ���b�#��H^9I`�TN�yO�F3|��Y.V^e[[��F��VW��&�� �9�&G+Ǘ�x|�^��&G7T�\U��五�>]�^��8m�m��4��n�&�DBN1*^B��0�ff&g�4ҭ�i:kG��Z<0�z�I��\��O� t�F�Ф����@�l-���~k��.�Wd,ll��4��׭���!���ݬ`e �Zm�e�l~]���9&���Oz1��b��UӦ�1Bf�Zfi��"�1"��VR��c+�O
#l�MB�뇿�%����ã�C�?l�eP]M�4����	������������!xpwwww�|�������S�kfM��^=����?�W𽳋7�V�ީ�^N���-lŷ?��G�\)Av>D�umt��^����l'T}N���PIq� �K�~U�� �s Zs²�� gۉ�}�a�<��|e�Њt���5IQ�1�mk�Ws ���&�H��(p.y��p_�>M�-]�����
EMǋU(�Mhj�M�3N��5�<f�)��u��ʹ��u�	�<^��(������^{GW׬���t�dE��{|��f�NM�q��-�!��,�+�9u���T���?���0&lL�0���)j+ 
�YQ���b骕�qs�(���P�w "�OU���d�����#c:BS�/@��g�xn���"���\����ʪ`��瀢���xN�+��ï�sdI Zw�k%�؃2�PG
�^�P��Tŭ�諌{2f;nt�.$T_�@��[쐑��7J"2��1���q����U��'���d"��CaE{��h��kZ�z�z�>��#y�����PϩB� "Lٯ88���,
�v���K+	z#��0�rm���ˍ[���_k�0��u�Q �j���I���mĭ�K��BXs����+谑uh�%ɖ��W�������}��r@��+v�	x���-�����7f��gM�$B�Z.Ŋڳ�j9V���1��ʨo��F;Ѯ��m�?ɷ�_���w[�뿀M���:7��f�3��vc�<G?���~w=5�N�\J���̦�j8�pb{���h?E��Y ��I��zΔa9����#ĭ�qg'�9B�~]'&(@��@��A˺�+t__7����0�&�فP� ���?��%��;�[I�!�W&x<���(��#`a����q���c9�,�!��Rv��
�c�LY��-(ɋ�w�vq9m�rS���mP^9#'�h͈�r����"�%��_��oI���6��,QI#OiK	<�^u���vQ�>���H�.=�dfpfB�j�uL�E86>���T��)�F:�vI�Z��|ߝ��	�9C�ъ���<0~o�ϋ��e�V3�����v��n�M0>w<S�>W�g��;�����T�DEF_5k�9�(Ia�D����`�L83SBz�蛎�[[�v�JЕJ{�0�݇�UR�U������*W�v�G�:������Gֳ7����c�N�O+(h�L��>�>n2)k%�'p�g<�lkh�~�!������W�Ԝ�����L�:q����m�l�v>ޮ,L-�����?vP���B�Zy���L���_�</��o`�6�܅e�:��g�9�6�ҭN��S��p#k��d�
B$k�*f�Vh�R&��*��E�S�ӬV�$nʎ��f��,eK��y�B#�:v�qz��
ًk���1:���7��|[cl���j2Ԇ����_��5����B~;�[ɛo�'2����_�w����ȅ�Q\
[A{�4:WZ�߅���8M�̭h��QT����0�B����[��~���.
��~ED�mm���}A����T(�jmm�=�9�g�ON�B������FM��!&��2T�#��	���v)�<=)|�x�����X��%��Қ����?ݻ|�xҧ����<@`��P���76��x�[_��R�V�Ij�;CU_�
q�AЏO�d�����X�Q���L]yy�_��dM�:8,	�l���Vs� ���f^��k���|��9Τ�X�(|<*���u�K�U qK��3��9�$_�gJ��l�;Tm����y��&���R[ֻQ��?eּzQE)Z���xf�~W�Ss���-(��� `܄�|���<�
ϲ~��>��)�~���P�P]���3h÷���0�w�pQV⧦A��&΃�]Ż�.��kpLK��	�,���&��^.��نj�>�v�Xt�hL����w7�ve]Z�Ԡ����_}�e�+Ȫ���ɪ���o`NJ�SN�θ���ڙbG� �W�0��Ql�H�`y|�\��>�?�vuW7O��.(а�:�'�lQYT�{b���Y��o7a��Ru��EZ��D9����gǍ����ɹk��yDو�z�qz�Ϧ/7�;�Ztx.��`�V�E����NX&�(���!��+�lٶ��^J����G錸��K�"FD NπgЛa_���2�׿�YEH��h�2�[�S/ʠ��B���4f-�4�;<�[H���u/`����]�3@~<�*0�/��l�SQkvz�E�M^�1:�I���I����TK����q�G1�C���3�j��-r�\8���I�^�v�t���aj���6�sd�\�+�t�]�{�_���nP��}��}Mr���mx��^N��K:z*6�8���e���g��3g��m��JS@Q
r�sdC�b�m�@��k:udCc6�ED��׌&y���d[�mB�6�d۹h?g8y��(ʞ�uߗUhA.��i�@��/��Kss}���€��7A7�5w��r��#����}n���磷���	�3�K�.Ol�`��t�z_���@����$
\��˺��i����]|!��_K�EL58�h.���d"w)��9� ���%��-�Rԫ�&��3��~��°���R*�R��I�
=�%Ksl���}���R����i��̒���]�3���)��)�M�͈W�7�o�?hTס2�(gcp�$vgf��L����g\>jf}5B�s,�n�{{yb�-�>�"3� �0~����5�P
C��d���7I�	����<^Rn9�:gq��:9T��(Ʃ�aj�7�����af:��~ ���+( "�1�h�R�m=��e�+��]���~m��\�ř�A��ǆ���0����[��������Dz���ŧΰ�I�˷��p����֨��Y�?��/��@*�u"��w2i��ްlkZAi�*c���J��]�8�uv�H���(�op7�+��7F(�@_��0o��Yb��&Zf�=��a�p�SR������w��}�ز��������ea�5Ɲ"�'�hH�L�1�䂞 �����||/��W}2���E�[�)������U�[��?��\����k��F9���oz^z��6��V�2J���k�ū��Z��	Or_ٞ��\���_yry7���@�� 2�p��ٷf�����M��.��;I3�OOφWp��b�����t�Ύi�+#DG�lB�.��>#�,��!����3xs�'R����6���35�˄9�Ä��T���o�=�������uk]��ET+\�,0��ѹ�Kj|���6�k�^��j�uBu=	�[?��o as�i���qI�Vm����������sV�Q�mf�-����lp�^�z��\H`T
�C���^r��.��Waͽ�ǹ�u����P������m#��2�����%WOl�Wm׬{.�K�F0��hrsC|
5�fy/��X�H�����Ρ3<SWl
�y��|��Օ���)�e�¾�Ɵ��N]���r\.t�W�U�L����
w4�5�S����BN��``BCo�m��\��j�D�_Dl�f!���~�� �Ib��'eR0J$�%BY��Ԃ'���(`�ӹ�"�Ш�gfwG�4:(����&\6���	�/��,����<�F���DS�=ꏳvc��g7QE���g�a�\E����?���$s߱�܎�͟����=6&�:�<����n��
Ɲ�iJ�>�f�}���j���y��"�CE�m�0f( 	>o���cЫ�iƪ)�e�m�Д��EH��=}��	c�e��^|�K��~sK���v�K(����n>*�4/�>�`�����EBw�D�c�ch$-@)�g�Mr�!e�_Ǳn���"WZ��w2�}x~�!�i�Ƥ��p-o�}��v?�9������Ǜ�3ऎ�<Rl��p�x�o�O6�~ȗ��h�w<���KO~>=��>�l�:]X���q�7�dw;����5<�^�O5�(W��C�B�����4c&6kY�^_)nb����,ϗ�3?�����ڠ���bn֗����&)��+��zfјl�ݲ7���SF���>�;zG�]Ɂ^o����́���/#B?]&;^i�>wS��ڠy',��w�D{LO[��/�/Wl~���ڴ��g=�������h%m��ǃ��H:�GD)Ք�#�cc��ޅi�ʾ����)�f}�.�J>���{p�~��̇?��>�Z}���/d���CCx�Pz�d�M�c��g2���8�,�|ALh�_z���a�4�U�Pо��w���1';/i-v,�>������� �Թ�gm�kpɺ1l[7Y@��������T���I�w������G!���a�ø����#�'��s3NqER�l�C*i�A3G���N?O&v3��_����՚��CIY���L1�y\	�@�󋢖�􋩮n]焦Vޯ�h/-Pڥ��6^�	vs��=Δч�3!���j�rP}D��J��I�� N�f���H��)�~Wv�1�J)���M��V�燠.��I1ɿϧ��Z�!�%�(�b�����7�v�/R�)l����l5>Ā�_9v�sw4��P�N�{_d��}$��U�it,aK�(Ֆ~��դ�����~+Yͺ���i��L'/=ꅅsҕn��Vo���%G)�q֏��
�BJX�ُ�P�QR���.>��چΖT��݁��X�ɔ �yh��ZgtS�zٷl4��I�SPʠD�/�	�Tc6^��cfx��G���6����f�_"���5���4��A� ��:y��-Z�R������'ᗐ�h~DO��H�i-�;�%�L��Z�����|��?���d"���X}Xq�rf�*��4�C~-Qߊ���e)���ˡu'�RD?<��C�<�i��^*�=�x'k1 �Z�1��*Ü~G�[OM�y�m�_�po9{��L��_<?����P�'�ꔆ��Eq�[j��#�Z�߂�!-��㈓[��K�{��AY��`g����6DWyrD]�-�N�N�PޗM��V�^=�Huw��u�E�*���c:`�:B^�jr_}���C�2d���� ����ji��͐#��J�����QY�X��22"�����(բe��ޑ�͊�Y��-������f�-�!�x��6�;�֚��"��k�������Mon��M4��&j4�����p5 ;2NFܲZ��H�\4�?w���N�Y�_
r ���@7ő�z��}(��F&��5+�Qi�8� �1� ���݈�B�D��:��h��@r�ۘ\Xg�	{5Vvǎ�Ը�_�]��1چ-ԯ>�g�Kpa/ �u�c���O�$6C�_"ɭ@G��d�(����`�{�W���]�iҲ�y$�`��3Mw�w�Bo�ٚ�c�ۗ�?�ient�`�-��l�;eD�M4���,  ���F�\6���6�A?H9heoY���n�,;��L����B�OeaV�o��Z�n�bu2X��t�<Gbd�&��ATbͣ"�ʢ�H��2���Q��Y��K�y`:��~9 ��-���׫$�C�X���PKo��Θ�y���,Ȅ|y�M+S�y���?���,�d u�U�N�5�����'���V�8 ���Ͷ�*�/}V�K�)(��\���V}k2r(���t	�� jZ����3'�tRey,
��"K ���b
i�c6�_��P�Q�S�!�ٞʕ��q��~������Y,/���"an�挰񃓱���fcd@�߉;�tE'���5qG6A]���3h3 3(I9d�1=;�{}����k�h�J��� ��[V���1#�t����:Ǿ�5�Sequ)����t��NR_QUT���ravfs�x�0
�!*QXD�i�M0DT;��ۧ�r�*�w@Ϟ+>���B�[�;���~@�C�q`����aG�U�af����p'�Y�i9����6YCW�\���W�0˫FOB����k�+�<N��44�q����E|[��žke�ԙ_�:��;�Bh����7kv��qgqmh�H3�{+W���`��R;N��3��o\3�Q&k�%���;Ȟ�NK��>�$�pZ���n6���+(���{d{������?��2�;�Æ$�j�1_��&��O��C�d>�ujGLSM�j*ݬQ�8��Y�9��V[�V�XA[{%E��C��7a�qʣ��{w���` �*_+>~ʃC��:�R�3����p�ם:s���
���� Lx�_;y�Z��_0w����!��iD2�^��g��Sɔ�qA�o`�Յ|��X;���+�*wq�����FR����j�����V��R]�6&�#{�<H'�Q�]T�+?H=Ρ�z��%P��EE�2�%VeL(l=���/@��V���s.�?Rb?��&C[���%��sw�C)�e�������NR�+::�|�6H�^����'�U*i�R��g��i�EAabzq��l4/�/����[J
��R�c�p���8����k���� Q������8�^�5�z�����`�Kx��"n'�sZFN\|wΟ'U�o TFy@z�;��Irq˭t�m��E=�}5�� �(�*T�hqe�(MRx84�P<��~�dqzH a�|?�\o�!�MM�׀��jt��~��9��m3
N�AJ�H�!�(�h�j����u!��:����Ry�J�V�(lq�#5@��nB�My��'B(��:��)�Kl�/x��f���Q��!aaMM����3N�zu���ɱ�Սu��w��K�qL�𹿔�E�~p����dnf������o�-�X���w���.f���j~���:=���n��.f0Xcw�ÛI�@�Z@q<���.q|\aQ�fi =M^F�8�����p8	�O�b�m�͉���3������p`�`���(S�d���d�������MfU[97k�!�/Rʣ@!ա������R���f�4������z�=��'�w=u�`�̉�0Re�BBD�seO�D�D�ʈ�g�Lb�_2�b���4)k���C֖c��-!�����E�>�uS�mT��O����w�S�V��>J�:9��([5�²���q¤�>�ag'���!��Y&�o���-b@>9�y�F>+�w�FzA��
��=������'�M��)dcgg��#<����}`�'P�&? �����ysr��H��7����,)�D��u%���,^�"��j .���]GP���ܔ}��
הM)`ǀ>�H��� e�S��b
c]3<���|hHyV�7E���r�0�ה�R�@��F���UD�ʟ��3�	��ϴ� ����K�����f!����Q
+9&��|�3䰑��4Bdwz	�W7C\^2��g%j&���TL�c؁J�{Ϣ�%Om�T�H�?Ū�$��ʴ��gf4���a�UUA>-�Δc�Y��E�}���_ �c��fi(�@7i��8�YVJ	S������Q��4k��~%���M\�Dd�	y�������J��KG�	"�8K
���J�=�b�=No��i�0dG*��j�b��\��iz91=�4�an�8K�|F��ٵ�d;X���,-݀M�)yXz*�Br��8^�N!'�(��Rt\���Px*��N�e��'�:�z f�͖��<�rh��(��k��⢍�j�7��z����g1ϫK�[W����0`���/�?�-��l{?Q�Z�.۞q]y&�X�B��g�A:ը�	�
��u�$����$(���R���`4Ɛ��ʤ5z48�������y�9�lvy=)����f�ަvmO��a=���<��Hʚ��	�H���|d_}1�-�)��Dw#�؞3�:0X�"k^�R�\ā*]����M��r�
�G��B�prpH�= �Y�bmE���9m���d�ഺ�06&�^X`���9�Cfn��F~?�k+/�r�͜�)�~�F�GD��}l+�U�~[��F��tԙ�
L�2p%�9�+C7��4�F%�^m0�<�ȃ��b�w���K�Ф�_of�6�twW�}���zDҖ[Q-+�a��X�Ex�s��au�^L���_�x!3�|q����:G9��]��FO! �*\�J�Mdzc,�	Q����J�bz���@4���o�I��N�u�k�e���^�������K:l���m}	M�}FО9�[�I����\n���9�����x���ʟ,j�Mx2���+g9�@��{#OҘ�W��d%��cG��8��R́@�}:�,,,SS��iU�R�`�p��%�8<a����T(D+��ə�3���+������؆��
1��U�5�+��Gl�67�X�GjI|'kΡT0�� ��Ѕ)n�v�Y�!�\"�R|L���(�lx���'�J9%�F�-�}KB���=��3������9؏?&�*7�77cy�* �\-��RUb��n��Q�Vӡ/j�/�[��m4_}D!jxj����Rƶ[��w	Uj��_���ɑx�r��HZ���OR1�U*�X�B���6�{v���7#I���'Yk�گ0x'��ur�������ܯ����ó<��&!(k��=�Y��F��L�����A�6"���8!Yc�0�2��%Gkz7�菦�2��ؙ������N�y$��yhqd�@�2����t�c�]��d���7@��d�q�%�3��)�0ǖ)�c���Wn�����y3�63��Țs���%8i��5���#������@����O���oj	��Wب.��@���@�vc-b4�I�9�/�XS� ��ѐ�\��O���]p�������VQWY�A�����`��n볯�nMX�M���>K��NS�A�*�#b@*�?%�)ֽ���I��y�m7��X\�$#^�	��!=}xM+K�\~��&�WU���+��-<���ѺjP�\�ͤ��5�馌q�X�I�J�=A4	t&�}^�S�I/ԡ��2{GprӍ��&!ֶ�,�o�����S;b�>P�����E(ݑo��|sU�ӫɸ��7��߉vX�������x���M�Q���P=�~t%��f��a�����H�f.�a^j�uF�漜�c�;:xp�!x�
d�#�w[��y[��l<!%�6TײW���e�ߑj ���<6��,�4��G��B��|��]`lT��9D�}m����@�3�%0,�Վ��:���Z1��P��.�]��bj���V>ǲ�̘�����L+-����<g��&��%��:4܂��=��?�}���h5Ĕ,��nX�������vfN�Vc#�ޚ����� A^���yW\2��	�&��85G���_>	;�O�n��;#c4���F�j�2�rHJ.e$g���hc�2&n���6�_/6��}�,^�9���;��R�p�.�{B���ExG�5����B��;�Fo��/%И����fA��9��ґ��wb��.�5�0��id㮍�#�8E=R}�k���`��hj����Kv>��UesgL.�_���U��p0��h[��#z��}M[@�G��@T�v�c�[깷LbO.r�/���+t���;6%�ӹ�4��i�_�ZD��9	`�B�^S=>z�����k����M�~V�"��s�)��ʋc�pi%EC�ϛ����ʮ�m������(<�� ١������g��(�X��b����t�R<|����n�ֵ[0��0�~�6	����1�	f�m�q
yo7g9�i�k|�K��,29�d����b`B?�{����`�=^}�c�Ң'&	� �S��{��*L$;��ք����CC���	x"�/[�B�9��қ��IQ�i��bdP=�ZY!�J�I�:?'N������_Ǘ	��?r�T��>.G+V���6�� �C.A��i�^�I�Ac�Uj��A�>ٱ��A� x�%��
a.�D�O�H7)������z�p�Wj�"CI�����y���1���\:Щ��"���[m�7�(Pʈ���e9���-�!E0�2�by3$s�	���߽�8��d�~6����N�2K3;@���
��H��1�����C�B�rM��blh��� �A���@V���Y"����ѻ�f��dI�)�QRn#�a�t��J�{f����	���C�곈�㖈%ѩL��	�U�P���g�����p��嗔H��a�i�7{$ȔH��7ܻ����x�EG��c�E�x�*�I�P�(��|E�#���m�,�#>̅�Å��*W��>u�ւ���HN��Ԟ� 7��B� �RżtL������K�g������.��VB���v����ڄm|� OC�R���v��c��`qU�F��"�p3
�j��%E]���XX��-�݆R$�dr@Q���4#�-�=�& =~�)�#�p��e��e� ^�،��9�h�n��~�rQ���&	n */�ݬ���gD�f�4�Z����(:�Nh�y/��]�ػz�T�x�#�?�։��B�)=���u�eт	��*rPfS�����O��W�JӐ}n���d�}�
_Z�5f��}F�Kh���ri1�#�a�'���rO���i\�fo?y%j�P��1�Ou���0��,�mMc�z�r:��蓜q�A�����.u�~^4�b.��. m����V����_t��4�饌��o`j�g���H��Ɍ^ZQ��%���0���iϒcN�]�i���+�\��-�xu�:4,�SS(} r�P%��8&������f�������hY�e��~�5F�����Z�5s���!���E���)f`[���7��_\$oaG�K7����+	���a��(%����7�ׄ�vo5�ds�>2�ӻV�k�'����cǽ��}�?djp�v[����w�(�o� v���1�oh���)�z�����*�- {e�=����o�d�}�0�y%d��LP��"�W|�1�w��c���p�M��������aW�L/%:O!�F��F5�;�*$;mE�+�A@/��'G��ȷ�`̎�k��ӷ��0���E��|a��c;�}��bFKj��������U��_=���G쫨$�yxC�'X�X@�ճAX�2���!�K�r��jŕk���t*��J��v!@����$����Eh������J#�#��s� Ӌ���tC�q2QHj�i��r�D���#ʖt|)�$�`[lLD�������EBȟ��4F%�<���P�ؽqJ�0{؛C��1QiO-�V0t�,C:j=�V{б-wm�/��60`���O�m���#��^D�{s�ǻCgapS�	}5�	���x�li�eJaY��G9d��[s�6�d]����@����+�AR�E5��(Y})�k�ڪ�=� '�[Z_��KS�"��:9_\H_lZ	Z���N����3I�t�đf����C�e�aa��ɼ�+�LQ�" �D��pؽ8?O�w��H�I��؍�t[|8����� �Ô��'UF��I�ٙai�4\<yY�"��ܥ��+�a	�
Bv�!�����]@\m�u-�R7S7Z$������H(9�u} �1���Y��k6F�Z:3p�Oo��(d���5p8p�}��1}��rtU���ߦN�'?�VK>CP���6�l]��)�b��꽥zb-�0{��idx9bjqaR�x��
����"oq�.�Tn�/Ϧ4@����d>����r��[v���T!P�R#V���&`��ʤ#Vϟ��*��\�X8��#-�r�)�"*g�ݲBNսe����f�KISQ+ý�������X��wP��M�,�,
[����c��s3�2$F�N1�ZwX��zzug���lW*mS�6�TL+��[Ȣ��ґS��v�����W� ZB�xs�Х +���@�r���#=�|�jHcOf�@?9%5]�5d�{��U��-�ts]�Fm�o�u�o����t���k����1;N�*�	Y\�%�MGy�f�:m�5c")f�2�I���孨�u#����d�1�s
.�|��N&9iW�N^ȫ��H'�gP�w�_Ӵ2��.����p��+�oH�&�����\t��5)';>�ds].����J�"�4|~|�:ғ#���E/���4ؠ:؊Ƃĺ�t�*�a5��\$�X�&E��|~����#lS_��ŧ$�(�Ç����t(tNQzA1�\in�uAZVJ��!��U���m���I�_��Y3� ��u?�Ќ��fn r�K���)�z�C*�p�̢�W���ڡ�NcN�	��"f�I�x/�(ϛ��#~kVJc����<�H(��p5��v��R�VN�h�eF���6����2E�dh�RR�O�Y*�\�@�H�S��E���
�UH��ז��<��,���1(~G�T'�T�����/A����#���3}��.�=Y.�#;����[�b֡�����l��m���t��:�QձmI�X�t��� ���+4�!S�s;@�άؼx+�Ҡ9�5���㔫+~cr���YB�{�DE���w���k��q�>�w����;��N��}�g1��"����L����<��0�fN�ίH��_������:��wtUP�"����'�[E���9�Y��в���uc���rd��)p��������]+��RR��������:�5�J�?"����M�1ܢ��f;�l�֥(5�G$?�g��P8���`hiy���U�hphU_�k1�>�WfGv{���`f4�\�\��
�:�E�/��rU�����eQX�ڼΌ��"�>���^�*����J����	���8eͣ�9�+�f'��U$ UW�/L�<�R\ٍ0���1O�W�0'h:oTQbn����;�%�q9d��]o��ZƘ��|BSwkۍT�����@�l*�	�\0��������:��O6ߦo�8�+�̐����͙�N3r--J/��qw.;gb�b�o�J�CG}����*�lC�t��MA�u!B�"�N���^�pSƪ�_����v�a�������ߡ�B8���#����Sb��B��>;Y{��l�O3\������� y�=���v�4���?2TWV�b��Q4@��&�ҋ��k�������S/�v(�{�n�Փm�u��r�/5����wԵ'0=�@�}ٖv����wO[
/��.�?I�ߛY�7	�L���uH���f�}Ip����2�2��zt�g��V���V��I�Ƿ�~3��͝@��6Q~B2$����Z��������|���;P��G|��>ʨH��.�P��xT�a�]}3�dL�ѿ���xI����O��Q����CRe{p�:�I:t$��?��{~k�G�&(/�6c��t��K-)È:��zX*���W�o�
i:�7�ћ�����ջ*��[1ؓ���|���:��>:��54D�?��3-�n@"ۗOI߄�S�RT�ʅ9P��*�R�YC{Mb�h���c��Q:�|BH�y��+e����� �8J|�&���m�~
��2�F�G]���7��3�}RP���q�"H��|��������uv�f_DI���^�Q:�;T����$�gv�Ǖ�n[�����b��2q�����1֑^c��&!hn���km�4��t�'� {��W2��3+ǝ���+�W�ٓ-Z�`B'�w���ߜ�X�%M�Y'�n��!׆�:��G�f�v�ߨ�I���EE���Gp9h%��wn��P���)�����%��\����*mCε��8�w�?�P�0���� ��
6x�c��fn���G�|�r�r���_$-Ѣ��*����k�jwc�������E��+��7�ʭ}�*����eR��&�q@-���{��d⟥%�_!��s����ݢ�i��*(n�S��������6yN@3��Q�<-��ؗ|^q�/��է�z'�-:�&��.q���l9���_����=��b��bG�s^����^��	B��z=T�yl�����~��<��b��/�_�
:,���K��M ��j�z~��ޗ@o��~�s��:���תM��g�>��c�	J��`�=I�?�|B��dddY/9.�B�3��t�@$A�����8�a�;���͹��N�V{�ۢ�vk��S3���B�3���Jf:x��ݦ�3%!M\�d��q�_W�= ��@d�d2���
n��Z�d�eΠCkR[�>�ne�b�6���u���_�6��O\�z�G�h5̆�<S�ͽy����� ��y<�X��庡����Y�l�w�R$k�*ⵐ)����;�:F�t���T�%!I5�wgT|���Q�u�����"��S�e��^�"���Ne�.R L��1D���VKq"������L��$��Jk����ٯ��$d̾=F/�<�ˑ��_�%L��5VRs�~��`�R0%E��<���*q�_$Y&܁:F��*�҆/2T�����/!;g/}u�g��:�9E�k+��L������MEZ՜%����+Z�������ft�.Õ�+�ͼ�� �V=���������d>O.�35oe.��"�Z�#tp�؋��t�/W�{Z-��v�����q�{�@_��#�P��)q!L��_|
a��N2&��>~����~���o+V�^�N@d���Ɠ��2�y�܈(ފ^$8E��01육���<����S�ʏ�%��լw�NG����̐������P�ǐ�~���~�#x��4������<OP���t�~�r��~���)Em츪�9����`�4�j�r�X�;�T�=8��&"8�.�Arz�S�y�B�P"'[1�O�85��1��o���)H�E�Q�X���V�:���֚�}Wc�^U�/�7D�G73���:�#P��o^��>1x�>+�wH	�Û�+לr��
�r�P��+V��}��EF�y��8-]N�B�^f/��_A{�&���mCt�U%�>�5�[�������k�D�Q^ʭ�r�O�<ai��\:����]
�w;\�����-��U�E������j
P��zO�{�\��$f04.�����d])x�4�Bc�E#��������
�*wH�"�7M/�5�"��NN8�s���������5MBoo�y]�߄�.Rz�5@���B���0��+��]s���>���'�4�VꮾT����3��p@`�t���r��^�X �Dy\�9�ov�
���8\��\5+''%����z~A�۷$�e���0�<)s{B������MaN�+xV�T������8���s�����1tE�!	��m�1!-�����a����C y�<�"�$%��$�GVVY�|�29r��
ZS�ӳ���ޫ�<>$X���a7i�i���f�������r�� �r�6�1���yD�-}�W�@�>�'�O�QV�eNpc��Y2g�џA�4ƌtf�ġW&�[rDK�K�[u}����Y�M�&I�1�z�u������ =�b�/�76v���c��=HU���V�b���(���"�V�3�u@ʾ"��e�u�l2�*���K�a$3J4�	����?�`#d�,�����'�gj�	��*D���?~˫�	פvԛ����F�� �/P�#�
Z͔�r�E��-it��G��IB���Ǻ�xU±A	w¥t��rl}�������B�^�,�:͍�q!���̧� {F �*K�*ƨ�x����򸰹� ���_�}7��^�I �~s�?�ۺ9�	?q��f�?�,$�v"W��B��r�2I�2?c+�KZ��Ʒ��RDH�������0d��\yon�ŒV�߭b~l�����T���	[�h����FE��e����-"c�	yp���I�𵚰�qN�bvЗ$`��d謍0b������0�P��8*�
��*4�h����]'���Z�Wo����s��2s�?n��}���>����#�Խ��+�
��j7��Z0L��-���Q��7� rF�|���+�˥� � k �P�P,�}��׻J&O)��܂3l_I�FbJ`�#O9/��P�Q��a�L���M�j��޼���6Q��h�gϯE��O��7�D �'3��n��lY�>K��b���BkUnܞ�'�w�<]���}=6���
�f�n��[A�,
h��,�k�--��5r7����Qhi}u��<���Z{f�y�L& fR�T�0q���]����SX�7Է~Ξ'��Zd�1��1g�\��!���i^L�:S����Z=��]���>_3F�@{fCv�v�G@\V��,.++��E���#6vz=����OHR��)8"`Z��J��m��5��#&Xa�2�QAn&Y?�!�*ʧdw������:��,6i����nu8���{Ֆ�m�t�[�����:ٮe�n�:�Ʋ]�g���=�}_/_K��\��;��'�7��Y�hVhDy�}\.�(�]�tT��q�|��$�������-��~��DIƬL��+>=��/j9�r�DC���[e��$�ⷶp���.��'��.���aLDٌ?hLL�W1J��"���߿[�H���UWu$��9�h����:�"�����m����}�6J��O�2�2���ۊ<1"`V\�3.r�18T0[Z
���.7�/�~V�B\\
��-�T���5��N+?2=z�؅�%Em�iG��i]w�"��O �KI����z���V�*3}k����;���b����d�g��Z�8�<��W��:oV���,R_���~g����>Jc|�-�"��U�/�Yw�g}w�'�z�nk��u;fS�Bq��j1��S�����o(�]b���8x7�1i˹�3����;����.��f(`'��%H�yFx$COLr�m�?��4[� ܻJ��zi-2�G�{YC��hq̌褛~��{���3b���=<�`��Z�X�
6uHJh��$��ϊ�:��M�
�@n��J�|�ZF>N$�ߠ���֩�W�����߹���\Ϣ���U��ᭋ��"������(���^ʏl%�HD���(�P��J;�<�����~�7] ��Um��zwG��X'u(SyGLV����j��^H��T�vߝ�j%}{�V�ld9����	�)A&�8M��S�<o[[|����羜0��ƁB�"�Vp��ˡz�!}�U��cG�f0TX�bbG�_����X��$62���%��`�5��K�:�aҨ���5�Vh�8�hJ}� ����p����ee��U���517
Un���P�<.���"8��8��eutTJO�iR����0��K\�(�8&����Wc���"S�j��rs�z�ֵ��>A�_�Ȭ8K=�$$�NN��E�¹g��� .0�FUd^�<}Q=��ej0�)�W�v��[
oySMUgG=^�Jz}U�Fـ�v�aN%$�P�_����_!����_����H�{��+��E`I~�|���t�?	1�g�'�����<D�겾+�	7a.�=���0��D�NI�ڱ�,��gI�����C,'NA37�G�����P��le�� ΃_Ϝl����(R_H�c52��X��(��>ǉw"���[o�
܋�H��t
.�)
���Z�LU��ˤ}}yyM�D�U��]�X���o>�Y���9�6�RTD�U�.t���Ii�}�yQ]>ś+��5���H�(���h���?z��4VcmwW=q���p�P�� #'~s��<����[����W{�v�啓������;��ϡ�k.�N�R�4xH�K��X!�Csݸ�!�WR!����Ȏ�,L�TptX)W�i`�b����_�{���(������_r��[�{M��qe�J)�Q�7��[�E����cE��P B'	h=g�'��~t� �����8F�����n��3U��Q,H���&�E��v����8�u`��ִ��`�:��U��ڧ�-Um0$X�����[��E�h���u�R�d�(ʣ<���]�m��6i���ῄ��a�yS�&x�4��y&�pc����'fi�4�f#��88~(j�z���e5�b��J�ά�Q@����־�h�$'�V�XHC;[�Y�����}A����Rĸ����%�P���A�Ya�k�4Q���
I��o�kd�df���LN�Z?#��5�M;N��B6��s�O&�-e��r��`%>����ؑ�Ƽ���fܼ��y�^���� kmPI�	7ߵ"h��Ryh-(i��Z�O�;D���C�Hb�K��!\iĄ� `RL�g�A�5�;(~�pw���	U/n}�&y�]��4�$n���ۖ<�Z�8.���Π%ږGS��!{E'�J�o��V�	
����GN�DHFK����z�b5q2eh2J�d�M@��,r�H�v�HqA��x�� M�=򤨫#��q�J��gqݎ���6�U>>1gV�~фH	��+7����u�80M�s
%X��}B^!Qn��K���r!����U�U� ��̫[�")�IE�/�m�v�:�?���+V����=LJ�DP@H���GD��4���H����c9�@�'8�1���1p����wZG�{��iEg3��
�
Sy�FdvR��w*$�T�K�VjM���͑?����.A�g\��C� ����8k���.�kC�â�߫A�������)§UUp����~��4W"�4�=��S�N���eL�*��Z���Y�FT�O*����	�Ƅ<2���F�i�+K���~��őTC�Ƞ�U"�M^��Ċ�}�C3�8j�;�n^M�U�]��Sx(N|�,�+9��/����}L�8�rw�N�@B���5uix�@r�:�>F{�R�d�B�7�l���Fr��}�y�X����_���0��
��:���ʹF��MCk�àN���1��]nM*�ɴϣ�Tp]9g�D�t��y�k"��z_ܽS�;;+�0�'��K^�OZ������O�xf,�t.-��Tj�_ꫭϲs�;�f����-�p��^Ƨ�� m�:[y>�pu�2��X�j�`�|G��"����ǌ����˔\'䦘p�A@��G���G�wZq�ʴ8Mb«$��[^HU7~�U:�<ʣ��	�9U4�]B�Z���%�3
�,�;��撛�w��^�������`��uD�y::�[iϮ���c�����q��|�w��&���^v������������Ę����'�^�(U�@�����
[�5�1ڽ�A	����[���>9�V&�.eF��6��4�����-�$A.VN���e��������{پ]��j7�����{��qsճ!/I�?�`Q�N���5������:C^�}���Ō�q�c�Be��o�����[���e녶�8_���;��o`s��6�4�=��ٛ��5Ez�RjV��P��PV��O��''�}���@B����4{���O6�A?߫�n�~�����8���Y�5VX�#������vu4��ZE�A��YhL٩f9��e�^a������=�D���:�����AJ����^Vv�>eFhВ����������+q9�����H��k��=��m�E� ��J{��ǉ�e_�t�+���֞��T��������ׇz�{�ZN��.����� Y+��щ	�l";��9j�����?y-rM?%ȍ�ͩY���_�<D�d������5f,��-[CE��C՝Y^�4�e�>���I�n��&\��
�Nہ�=��ӟ����Xǖ6w�o�VO˺P������I�Cq"+���AgP]I���G���������he�1�[:V��~��h��X])��z�7������]�U"�u'7�,��x��(�t��7�AE�kӰ���ػr���Pܛ���:O�ER���!�ocxX\�Jbu��u�m�?r2��w�/i������. NJ�p�ۑQ9���
�?���?릯z{��xFҏ�����:�.&s��-�!�!�,<�*S~�=�'����ǖ�fi(��-��C��l����;�d䳴��HG#�ٜ���~Jv����1Q�y��s�D�j�{O��!�FS;��%o}�I�Թ_��v��m��`�yW?�ݧ�ӗqo<�����W0n!���I?�XBɿ��EX\BSǳd9^���<�~ �O���!�i�vP�����fF_p�(��������~�z�S�������MRnn���P��%�ń+ ��4]%m��a��DG}��cףߛ'S�b��G<��&��F��>����֪ܿ
�=}6+8���E����Z�i�xŚe{3�c�D�V�d$12Д�I���RMF;�⼷7K�z|��Z�6���~w*(g+��]�/��aB��6\p�����}�Z�~�95(`��7��Y��r�f0�"�uܑ��F ���D�V�1�p�ҌB�"�93_�#T���.�S&º�rrF����_QE�4���=/��п�{�2��Pݕ�����^i�����~N�st��g}izT�?������_�*ف����b+/�e�����nߜ���7u� ҍ*���A�D�g�(��ˑ��[�k��U�Ģ���P���Ȧ@G�'�a���,v���W@�5�$�}GZ&��*X�����H�dx�7�����-x*����# ��<0O�0�d3��>����j���IS�A	���\���;A���M�x7��x
��u��|.ǷD�y�.��Et�b7�Ȧ��5/���K�n���_5�z��)+^_~�X�c���E�C����߲��(q�O�=��N�$2t�=�g���!��sN��N�`'�x��G^@̂��M��P>�XNC�T�ۯ&6|X�&U!&���-��V�S�v���qt��y�#���7R
�e�-�9m���L/�I��C6g�m��L�2�!�����ϑ���
�yk�Nb]� }��.j͑�έar�#WT�����S��\�����	����D5�	h�ޚ�7�F�e���������Xdp��ą��ur���-��r��Ru������<��&H�!��:��n�ˑ�ZY�~q��|9�p���uyw��2S�W3�)�w2��_N������Vt���̕++Ktq)J��������Nu�����m��&v�
��ĄR�j��R����tEdm�,���z��Xm�Gi���^�B?�U��۠kbi�w"���#�*�hҥ"�3^D>1��FﳂL������������@f,q(� 4@�g=�R>�6���ʹ�nT�OJ�?��w�3̥��|��'��%z��y����{���4j���������z��
Hf�L�����US4�	!(L9م=B�&I�I�����Y�l��i����1?�:���SN�u��������X�n�wxI�|����X���|�lY��ME���E
��h�H^��O��P�3�'ɀ�g'\(�����{����Fp�щ&0�y�@rr�q�5�S�S勜Ӑ�̌t1&�T�gq�d�x�MU��]f��v���Ȯ0T��+Zb �ݔ�G��+�8f|�X�
���@T~r%�s�Z!���Y���)�p�U>^S�ؓ�|qln[���k����l�T�����Z��m�J��;g�ܲ�; ��i�7�^������l��/B�h*�⁎��gNv���_XElQuc��N�z�;.˞��9"���D���ӳ�9N�.m7w��O����K���+s*�f�Q�~��v���m2��]mc�j���<3ڤR������֗E��Z�(�~�7���Av�c��,��#,#DN�8�|�d��2�r�ҔX)�=�τ��T�)�
�%�{I���8E�X�SM������*dz�K�ʫep��u��(N�J+Q.��5. /�*5�͋�:�䚳a���Z��6��H�z�" ��ڮ�a4Xi��nj�ے&�D��'ض���N?��ۭ�\#v��%mķI"�'?랚}�ķSK��b�O�!��'��'�
�S,	h�0�1��U4��!��bUo�,_~N-�LM�dāo]⌖��O��*��&B��6��)ҍ�K�O�ѓ/�54}��i���<D-!m���*.ϋ��PB�3�����V��Ĳ2x���L����<����� ) v�r;��l�ܷ�i�-�	�1ؠ��,v��!�t���^�'��^�~��-�|,�_Mh���f�s����vĚ���2���z$mC��د$D���m��^�<��Vt�B�А��8M	ER�:�?��7��,廿ki�;�IZ�A�kMt�5Ȣ*�A�{��)6� �w<��*���?!����>�3�yz3ab�+�=�:�(9�(C���z���Z��Ȑ G�����s6�tg��B����sbbZ������WH�
r��y�jE1�ܔ񦻭WB��,��ˎR;h����� G�l�d�`]EF�hw�զ�����w��̅�@v���"G.:sYBj������g��c��wo�"Nϟ<�5{ii�_T����p]a�HQMz�X��[�#��}w�m����V��>��+�o��#�:U>4{��?^��H<�]����G7����D4�#���&B�cڭU�T՞T^���/{��!��L'��]&͒G��}cB�Xg�m���os���+���6X���j��A_v98�\�yԶ�﫱ƻ'�bS�*W����0��O.�(��`5EО Ȧ��y��vh���BW~+U�E�E� �X�&��m&�#p��deb������D�"::��wgI��2MEf��o��^�ꐈƷ��,4�LM��b���iCU׾�:�$�2����#�H���hR\^N�YM��(���2�򁐑�]�oui�;N���z j��6D��\�дK[TY���>�u�09!%��_1.D}Ե��D���8��Jm�pݴ� �.��h���q����!P2<�;ʳ��m��L�,c�>R��3�T���y��z�I�&|�c[E��'s����$���I^η����e���n���{s6�}�c�.�LW�b�_�hkL��\������w�&��+8�IM/�U��Y��'��!K�C\SXG�ܒ�LJe|���	�S[�3� ��)����;�Ē<]7qnfY]z�UB}�LԼ\�<F� <�?���#��\�U�N��P�3C;X����%�E����� ���x�lhO����z�$\X>�_*��H���􉑺��9f&_߱@�^Z�e˒*�<���5�&�7~k�@��w�^s)�_�n}��dwh�����
�(&R���h5�����ZC���t�Tz��E�x_��C�j�J]\�d��i�Iٵ��˽� ]�����<P���pD��5V��~ń*�k'�{}����T���C^��yP8����j��Z\i�ޣ6+zltb��<�_��j����!�@�X���:�-_� �B���$�r�L��7�⫓�9Aϴ������Q��l�� ���H�Q�Qc��f���-U��(]�3K�������wn[�hʮ�T����O�䢫!rG��?�y�6����Ⴓ�z��Z�ImN�m�"���)bkN�=ө�ގ��%߃ۙ����k�s+����Kw��_trIn���L�fV���t��~���b��t�lI�,��9_b������ E���t:���_�mu+��p�vo(�cS��%*�D�Ţ����os��`w�}*{m���εo�������ػ�����CF���Χ�Y*�ݾ��͚Uf�h��>c_.Q���H>3�@�FB�y�7�a��^�
'FI+��̚y,EZ�>a�4�!5Eyd�5^X�+R�u����R�S�ٺ�n�.��ĸ��.��S��n@b���c(�ݝ�����k\=��|���m��M1.�����o�[�<�˜4st�nS�N�DWq��?���&wg;)W���
9�G�$o�2�)�[�s�z������_�����;y@��0�ߐ�W'��g�;?O�-߆��D�m�m�X�]�s�B��U��\�/G0�,�&���,�G�.ؾ�L?�N_��nלs7X�4d��h�Jp������v�7?>�ґ@4�����&��g��n��7X֟�}��X-��F�><�V�\�:��4D�/xD�?��2�vIg����X哴����������G�z@����Om�l�YM#6���)�%<��e�7���m��i�L�n��\2�;l�
���#����h�� ��E��*��3�X��3e
�<|�q*ѥ������"��F�D#��4�h�p��O0O�Ln��mVf���R��[J��e��U	=}Q|����?z�i9������/�<l�8�����`�o� j��OK=
�C~��gÞgC��$�2U��l�8H�/�����ܮ9+=\��~�V�zMv���4�����D�v)�]���j���Nx����)��[�3^�P,��`�X����
���Π���"E�I�Wq�Ƣmf���$	i���AW�]y�#&��<3�.;�'8`RgTE=����3U�"ijx<n���M�E�l�7�\2��&�dƒ�qV򓟞�u�d��n�Ada?,�����~s_S��Foӭ��V���D2}����p�:�W���%�[�I��B��Y
j��E.G�GγVF���慭�`���u��Q�M,2��C�Da�l�e+F�L�ax-m��B��D�cd��m��f�yS0���`�������3�c���F:���J��/��a!J��{';�T�g�ͧE�ǅԛ5��h�0������D�WM���/1���H;%�99F��#�1��i�E֩P҉sͪ��=G���y�����W��W����A�sQ2�����QO�vS�Qn�Ď��X�H����'F`Uf�����PuX����L3�T[*�m:�����+ȣ9ȳ��ƾ�˻������l�\�����#�d=W����.�5_���M�#u��9�����"hGr��C.���s������ZTN�>�x� �l]Qs�m�mv����؁�NU" �DN�x'�Q�#��>c7/`��%ϲ| s���^o�e���.͞b���n�~�ӧ��8�4�����<e����|^��1�qe�?�}x�qi!$�ř��Fa^��6,�p�Y�K9"w��Hĕh��h�l@��Ӏ�����&�Ͼ;�䙗n=�q�����ſN-��>� f���g�xv�>>옷�4�>u-:>����:�o7�Pj|��Zr�(�:Ak�F��Ks�[�ц��0kk�����^�&���V^�¿ƖG̫�Jw�Š�y~� 5����N�\wZT�g4\�[���!��#�\n���;AFF�賧��w�,��[��@74�뚷�>��IKۭ���tO[lI��Tǝ���:q��i��)�B��y�L��-F�.���>1Q����Ԉ�3#q���(�\��ȷ��k��:�t��+�l2H1�r��R��^�
=R���p.�>*�P��'4M�'3b�
�b��O�����{�+�	����w�f����� ��(�ն�f���Wh�9:�s!R���o����(P(���"�C��˸
��ܢ��Ew[�v�ao��Y�e�ϣ��G'�]�tvÑ�#?�[�1n1�]DEvr���c�:q����ӞRX�1��u��sy���͵1��7�	��!K?�\_��s�_s)�C��HK��x�am�{-sYZF|���K�Q��P�ӌ�����e����w`�Ӊ�_oF����@�և�"��8��^�-ϭ���5�(�t��Ɵ���J��ZT��a�ic�xaM�0�����r������h����	b�O�ubIb�S���.C�b�Ȅ}����?��!"e��� �
�W��,J'v��ȷd��Q�P�ڎސ�🪳��.V�Q�>,�BBh�'F��6��vձ������	�J��rB�Sgjk��G�����sE,}c��KKЃ��w�$�,�ϕ�/טBcJ��ٰ8Z��4V����n �ko��|l:Xp<غ�A�O摲��/�˕M8�e���s�6������<��b���^�����~"S�t�Y�;[:m�"�k�&���&����i����7E����,u�jci��R^�@��1ԗ��݇'���h��Pģ�{�M�+(($��$*(�S�k�n�ؓe�ř��"C0�X�<�D�S��������l�z`HV�+xZ�����x�LA)�j%���휖ǖ�٥�4��.z�Ƨ(/T�R�j��򈜄E�Y���c�YT8��:����''g3��Ȫ��a�����A��������~TM1���-�E�{���^T��R���"ɻ��2�5���v� D+���X
dlt��~I��\���G��lX�O��
���� thT�]��q�L�b�c��C�fF������{amEIf#��tY���>�|A����YT}(���7_@��H߬�)T�(^Ԙyi�	��ql��n�T����Z�8A��Q�f�&�%DEe�h�B��\��j ��ѳ��%�=�Avq||?��W�#1!��D+S��wĠ1e>�ķX��˹�>F�H���2K��W`��> �Vy���i��~��Dk��yM~�� :nx/ٹ}�IZ[����>�p�C<��Y/������2����j��K�ć����zR����-f:���+��F�,?�%"�F��Đ�!D�r�E���X��r�j���'�����Z�-�Z���	�͟X�E��8���.P{  b��Lc�/���NL��U&�����}ӊSN�e�䶚�\T� {U��H�v�A3=��\�4�JgΨB�9$�����/4��*M��#
m�a�{<���,�Xt�s�??#��2��0e�;�����A�� ���v䢳iw~ <���PT���Q������j��J���.�6sFc�i�_��W
�x���y��p�d	�C# e�7O3_�D�
jx���OmmU�%z�CE�LEu��Y���z���Z�����5����(�������=�m������'h�B_�a���*���f�b��ʔ�4�c��R�j���	D�o	��KV�о�Up��m/"Gpu�R����>�8Y��l�����e�"@��9dg�m��j ��\����9@��i��N�Kq��8w�IQA1~����q���������V22��dh�HC���G�1=��!Q�q�͟���KTS������#'Q㇋���"^�mI�>�+��6I���t����g�Ic�es
jC*��`���n��K����u�u��o���YB���2V���� �<%g��g�����ky���ͥ.FUl�U࿿e�с�a�`�&*9�q�2pB�cBd68 �X��B�UX;�S�u_�53��"W �鬍�4�f�����Nc����(3��[şO��0��BJ5�]\�a��X��R���ʸ�m��֢��A�ե��m���g��)v^A�ju
Bdt�o��8��k�N�[�.nnR;D<��̣WD@�$S��F�>P�K��ɦqb�
�f�?��iE���
-�\|�Q��e�XF�i�����'��ьY�Ɓ^�Q�8��.��P���*�5�N����W���WA��l��B���|�q�.:B��Γp��+�M�#�l���C�?U�;��W�3I�	���4�?����zL���Ա�}!���Hy��Ji����"�Yl���C��s/N�'��)kJO�-�#�a@�,Z��L%OĐqM�?9%ZīZ�H\�(v�Q| $,�@����R.�`��PRC���.�����=ZM�\1t6�� Ǵ� �amь#��X'�{8+n落Pm�[����	��	���j]GBF��+��4�p!4�U�_��̊�zw���8�r�c%61}+ɏ�+�c�*(𸂓�`�����K��R�H6
�XȮu�;L�@4&�2N��rM���7�>�gJ4��BKf��Q��<�On׳v�^�ߜ��)ѯ�
h�0�3;?:(����#��jm�+�9�dU!����ه�-̪b��6՞~���cn���e��E�lq��2��ZR�Ѝ[0Q�^"�m:gR���lE
��{�RI�����G��&���%��X4W�P�.�S��~�ѪK|�>��8�#gPgJ��<y�j���� 
�+�33��v�!ZLA!~�b�kvp�]���pL�.���e�$J�����ȵ �r�����Eq�;6v;��t��Y����,%�l� �u��Қ����V��FMb��r�t���'J;)D�1:]��_����:�m*ɳD<�����et(�~��*%�Ki�F{5�b�(�"�Ea$_���*�o1�͔TN|���
=�h���D�p�3�l��4/�a5�/�|��,��rz7v�4UOú�jv�ȥМ���0�zn�,l�t���!T2=P*G��9��~?��0�.T藬��j��7�gSL}l�D6���N�`Q�映�y�N����3~1쟜Y��6�o�^����3,w�}��عP�-w$J1��'�>�3�������������Z~GA���(� �w��22��c��d-��OZ2�������2�qHe8�%>�n4�^�l���MN�����F��Gp���''%3��Ζk�(��b����ȣ
��"D4ڴc�E?���Cb�ndR��fYCK��a"�q��%p:�0!F�a$F�e���h3\ݙ�Ç5��E�S>mt�O�K>Ve�����ݞ���n��1�!<�R��'unL^-��'I TN��ߧ+�ì���ZA�4^��q׍��󔚰.�*?���,�i�/ 3���Ts��2����5)1�\�vҒ�md�"(*�;D_�q@j&>��)��så���<<#��R[	��V�%�v Ќ鱷����u����2��1��2,4�V�`����b�n���`�I������ʴp��y<Dl	I	���.9�8I��W1��������W�m����>PP��f[j!�_�=/ȳ��ڲt^�\E�iK�P+n�߿5�u^�|�s)��&�8���L�D4~�Z�� ��4��As�L߮Rt|;���ɴ�n�h�=�)�/���(Z��3�o^S ޽
٪�V��[l;.���ۿt�	���ŧu���2�ۙ�hŰ������_��|s�
����g9!�X�_%�;��Ik}�S_����ޭ���O�b���{r��p��h�(�QN��D����>r�V3�6��#�Dc>5.�m������Of&�9ޖ�R�gk]a�a��Y�����hr�xxDq���űlV4=�w����%���u1n���kǧ�;&$]������B���r�c%����߾Y���|7t�}r?�_��%D^�
�}�
 =��>���A�Q��V�s��/��/����4�u��ԩe��I6VE�m=�:{֣��Xq^]n&��K�h�rR�{=�65�T�>����UX��L��$�g�
��S�� w��e�bmaг�vAB��}Y��-4�;�,_i8^~��D�����e��a��v�L[�jK�,�4_�y�GB�����3;�㜨�2U��l�t���/
��":������l��4Ȃ<5�:_�>���x�v���Z)�L��;O�|@m��Z�yѡ��qa�]�Ly�س����]�����y�I!���r������Q����;�6[����_i�0]r1�9};��e�ݻ'۱m<&�6%���ٟ'�@����Ş�T��SO�5�?�����t{�p�<S�v_4�Ob�u�e�p��s�浺��}�1N���w�/�xru? ���;��w���.�}�&�>���w���"�;{���r�K�����G��[��;u�����f�J��KDo��[_��f�*ӞF�qJ@e���U�ٵ�{��\�ϥ���L*�ț�5�	�!ε�2/���ӭ�Q/��F<�c�6"9������1"��"�PF�4v�4F#����9��.����z�Ͳ���kx���2EV�5�5v�fY��9]��X���������Z�D���������v�d�#��n�����g)K��~�_�����¤H�4pmԥh�g�X�+0��5��AH��3�Z�7��i;��Y�$ J��JԜ������y�rI#�l}�o��R\����8&�t�t�m;������ ᔌ�Q�>��ҞNE�^�H""���(�w/<<��[t%��SSK��.XԙF���߀o�e�/o������i�����:%8_��8t�9���Mw>��4vb���Ӗ_ׁ��pQ~�k~>KՅE{�����Ph�I���ڗF��7Ѵ4�琯	߹��c���N�>b�j�~V}����,m��?Q1��(Ҭ�D���XH¬�l�f�P�7��/�p2��Ӡ�>�i|��9k�z>��{���G�
T+[�ݭ��D�׉|=�5���9�=���8���7�.���&�(	�.X�ת���G%G��a<N�f�<���7���=��l�X�=���R�&F�\�Ph[)W�{�O.%
�Q���n��"KV�ro��ַ���@���2c=oO��A�G��3�����r{^<���:�_?�Q�h�F�?= �lAe�?��l���G�aɫ�Ia- ���[��k�dS�j��nF�1���W�N��^�~��m���������5��8b䶽�?�Yk�����'�M�n��bMcĉpq�8����\S��A)�['�SƷ��}���Jjr�FEc�k��$�Z��޳�Ve��nQ}�҇[��w�:)�G��d���Q����[��i�'�_8
:P��՘;.��.6��ڛ����\26�Y�7�hG����@!�~�`a��}	��E���_�L�#�dg�!ù���29NeVS:��Ebݼ=u|�uT�f���`&f�w<hd�Z��4#�lw���H\����ڳ��Q�������cbڟ	�[�y�^���R���)��î̓�@[���ս��p3tg��'��\���'��V]_tA+�ռ��̚(�!�wK����7u�uL;͗�g�0�{e�� /����J ���(D���i����(�Č+ׂ�'|����H�ᮄ����p�(?#���׶��:����f/*�� ��>z�|�|���y�9",mW-��]��b|u:���F����^u��`��;H�`zPQ�[�:"�K*K>;�!;��_���-��6&�g�[ʐ011�ǰ�G yj�a*|)M��ڀ,��,��Ǹ�0LE�t�X���EҊo<�6$v�<�zQ8�i�l��9�%�w��Z���fuJ)|j�&NYr��*u��%@G5��0r'w�8?ry]�z��h ��B���h�d�pD�j4��g��`�;���\��0o�Y)
5�l���<CeW�����8͊l�"�z�?&��(�>�5�C�F�V<X.?���Y����ew\v�p]z�~�3�����P����:`iե0w*��Vyں֐�~ȍvz��]���qo5Ż n?�������u��!�����=O	�/�{�Y�;ޫ4h
-6�7yd���$���f�N�D�����G��u P���W��\����Ի�}q&^
ڌ����?�S����G��SW�0�� ��YC�\�i��^��qO36�C��Z�qCkPL󔛃!>O�jf ���|`c��Z8��e{" r8����F-a:�u�8�oΆ@���+#L�~�d�ҩ��V�@�2 Z\i��ЛC�ˢsY�JSc�x�oN���!�@��K�L.��ʒE6�'�΢�ƺj����ݬ�C��˫�F�t{����<E�&�}ا)��K-#_�X��Ìff|܇V�l�\d3��!�\��#_b����,%�̈́�+EZ�5�rx�Ӑjt=a�(����7�������4e�r�*�(
]���R�иZnPD:�)����e\8>��07뒱�A�ϔr�"���\��hk��~^h ���<�Hw<���>^-��)9c������L�����'�e�;�J�k�T�e��	���p�n�d��x�y;py`6&���1XD�NР��ҵ���]������
׹Q�c�u�|�rJL��������1K.�yH�S,�-������z���7{������H11�8��a�]������q��r�t@J1���m��β�t_Lb�B��*O&��G���Vh t��6'L7�K�<#Qr�����:����%'ǅ&f=X�9�髾G���\!+�Cy�pm�ks�� �<˴�А|-X�cvq>A^ii­=�t)Y��������sW66���8S�5:f��#��C��Q�v,�!Iӥ���q��\j�J�]�s"��Q��t�J�:7e��$���w����I��qS���sMxF�Np�{DCl`�-^+�j8�c�p���7S/]�y8�3����S���8)�(�o�.F�(�Xse���A���>5g�$����:��T�������n�G�Y�W)�d�΢�`���b֟�����J)����BN;��l�A�9�F��/��)��앁�y���S�����;������׏��j3��ĵ\2�9�(���@�=���t���u]�xb�����m۞ض���ļ�Ķm3o������k�^�{u��v��ǸG��YoEj-�,�O���m?�L�m����>(1�H�.���-2pɒ�tx����[8�I�k�H�PH8ٿl��fs���Map����+P�G���uFiw���`�ɵ�)}&D��M�[����zO�Äz>W6>!Aʯ�e���l�>v���r�Q�X	�H�J-�,�ˁҿ��6��3Tcک��X W�L�H�"���,V���}�	~��}�;�A������.gL_�$L�kK/���g��8'�9���*���cI'�7������.2#��z �o�N�t�y-$��b^��%��k�s�����	>t�=��S3P�+��r��U��Dl�\�d�O4<�޽% ����q����?�Z�]����&Ъk-�G0�q��C/��H��d������W�c��;����t��e�����v��
K�\4h:�℄0���H/��%v��e�V�������po8�B�����S�5�����T��V>)�4�چ��K$�2�R�[k�^�֦�HE�nq����M0�8?�d��9�A}L�R*�=-��֫���q�~U߯e>���_���٪{�_bX�kc��HD�[�;GE�xC�����%��ZMN�iPi�x�}�j�����k7����n\\r.�ԖlJ���5R����e�? 
�!��Բ��p�+ҸٍЪ+�J�)����۹Gl�Id����.IH�{��C�����1Li�L�xfV�H�� XA/��*ZAa�&����ёp�E��}�!o��f~s�o�.�v��'���"u\T�;�7$h$���Ԓ��$�i�4��7�4�|��von��+��&�D"S(�RU�Q���/Y��?��"Ъ	8`��O��N9�-W���ܮ��a���Z��N�1����"\Pf0�����P�,����tU�U�U��2��4#�W>ym��G�GS;L���/�Veͽs����N5J�A�l=|F��[h����l�Z/�N`�)�d=I�Dc���=�Z�5[���K֚��^�ǖ��<�[Qr��3tb�I���pM�b�n�*N5A�ISS� �I��"ؠ)�hD>^���\M�9��X�_K��z�Z��3(;�9��AX$�1ܭE���3�s�Y"��{1=`O��]���'Q�C�ґ�"���bT5u��_��H<a/8�d�o]=�� O��{�����O���1riӍ.M��o�2J\ .Cxݗ�r����tz�r��|�Edm,�vC�ē�
c�w_��z�H�^�,�\ȷ�N�+�hhڼ؜v�pzZ�r�EUb��*�E�*���	?��9�-��t�V�)W.��D�o ��r�mp�@$7���w=�
xD1���/X�\�+g#Gn�I@���ĭ��.����_��㜯i?�'[{7:�N��Tq����Ӽ��[���H �Av����g)��-a��,��V��)8��|��y}f����ԁ�2�LT%��A ���3���	��E�}9��e1�4�$�d& ,�&��T6I����>�Z�ȍah����z[W��r���ףʭ!��D�P`|BpiN�,���σ��n��'-K�82�-���	v��0'E��:�@*���F!{I�5�t{��Ԅb����ְ&���[��d]��ɘ������}e?�v���F��ځ<uM��D�:F��VU*��E‬��������0(�B7L<,���.��3�`����`��k�D�Y�C�]zx���G<(	H�,����`R���tm?�5h�*�SGe���kQ8,�t�� �\Rd�.�b�A���,L(R�^lH}�M�~[��e)t��'?�T�n�Ь�]�&r��њ�6�WTD �}���N�*g���Ά�b<�Y�h��`xxR5� ����%yw�ErnS��Տ�h��IWF}N��i&�V�!1f�̘n��M�X�IpM:��������`�pbM�d50ɤ1����&�{��//^4��ǻ����<��id�=�Ny0F[���D+�;:L�Ce"i�[�)����2�+)��$J�(� W[4�������:2݅� ����7@��LdIϰ<�����Y��7�h��LY�Q�&��Ux]v=�x/[Ċ�_���*��	Wn���u�9��9�i"���Y�Jʪ6��G�dk�+Ѱ���`\X�2,7��<@��YI�0Z9Ms��!?)�VC�WKWD�n�B\�G��3?Z�mc2l�jc���K���KʝH�2M�����L [[�.��]MG�1��f_��lR4%����~/�����IIQ5�I�y��js{��ʁu�5��6$ZWQ�����2�00n��x�ų�󝓭aw�@��lo�ο
��L����*�Ag�1nQ�?�#��� �d�#��֏�g�y��X�g��F����ㄔ�����L�H��R-iEZ\��� {ү�"�_��܆y�Y���
1vI�r��!@0�(ϙd&#;W��E@��M�Bs�R�]e�f����m��-���O,y�'	�\�G�M��d�<�Vsj*؊��֖�K�������~���a-Wä����3+I��G�����_�MF�O�{��[p'凡��	4hiM�}�q��Y��9�=����t�a�R{G���N
�y���r�65Z��L]�N&��g����	^u<��\�DM�~�[�z��F���q���~�W�nv[C3���R��I`K�ggc�9Z�D�m>��[��s�g\{�8k�9!*}{���l�b`0���+1I%⻏����X�k�ɺ�H	�J�����ERF��?={9�*k&N�yd*����_	��U�����Ԕ4��I��x`�g�Y���`WeY&�Eܡ:=�鎜-*�ޗi��A��3��ZTD9�xP�t>�ʝ��0>��٣C���{���G�px���E���)�bDA��. �n���-�wWt3�%@���oW��Q]x��	;�u��)����1��Va���]��7;��D�� "Ǎ?+�=-���2i����K��^ۗ��OxY�7gD��e
#G�P�^���_ۡc��,���;C�2���
9����2G������٧qڙ� ���������'�Sk듫K��ɹ�9�Q��
��T��!0,����!Ek�}_��z�/���J��ϠNMg�+��p��+���p���ey[�d��+�[`Bu���,Ap�a�7c�˾��M��ݖg2\�+{'&cʄZJ��0�f�U�G4@���tm��aL�{ހ�s1�1��̊�s�]{�zk�
H#ff�D�N�b���h��%�)�Bf
���0��tzϠ���>�E�A��2d�����%��쁾d^��J���,vpw&��$�8��ѓFx��yG�`�0��Q�<ʚr�R���""�����U���%�Pm��K��ܪ��p��}޼�6����/�Q3z�rgO��f��(��u�6�֮�,��p [�1uH�>�L�f�#��)��
Y�}�(�Ɉ 8����Lu����r���գ=��(�k��װx�y#G�2�%>�g⍺�ĊMD3�������U �D��Tf�F�7�q��������)6w���3�U��{������O#����"����m��W�e#ż�Gs�m������|�����,&�=ڕ���ཞ�KT^߲T�V�ۢ��_��(���,��l�!�~UI?��m�7^v�M�,M��nI�|����ڰAq|,;ˉX�p���w���'MF�}�et�H�0|f`��C����\�1@�
Y!߬;�߄&he7ߢ�'g��n/��j@���7.qK�M��;6�A����o���K������֑<~QOu��ם{��#�[}��$?���X^ˏ�,$���_���ui��!�/8S�v����q� X�X|#oJ�n�?�%�)���>b��SfM�l~����%���6�PM0��� �1?��zC�ؒ.HN��E[Ogj�}<�n.��.w��Q�k�[=�6s�ߴ�~kx�]&���H`�+ug
��	��#A�!j̎��,o� R ���o������kr~�p@��
X�R����T]?ŖSWg�l7���w��}m�#� x���=��/�_
(���S�����{"������4��1Ĭ�[�F����y�L�P"�\2�7b��G�Ǥ�K�)�YH��4�T7'\M1��<�0
����y������6h�����?�l5E�F$�g�{���ܔ��!N	�J�x&"zFn^��a��q�L@;���4^�����`���hݒr��A�֖(4�e�J���Q{iv��X*q��pآ&�j9��#�����|vZ��*U^�R��.�H QvSI�Nȉ�TSXP��>���^��s��m
����h��#��D�2���I�x�"A�'ƎCU��=G����_��F�ٿ8W�X(�
�(T'�)�e��HA�])]jfU�?{O�>5���H;�J%��P��/9��bE�οs<����U8_�˟vb�#�G��N��C�^'{���)�n�
&^E"�oW��7��w�D�Q��M�`�6�"R�j�d�o�NCcF����ԩ��)�����4���{繭���Ʋ��xl�{DN'PH8�`���a��<���/vC|ᡠL 3כ��ڴpO���HB�'��ң���l9�����ħ�)tpu1�rs\b����N�O2Sa���3S��y���Z���?F��"e�c��8gu弍�ɣ�fW及�w�9�OE"�Na�]�K��[�e�^�츰�w�Z�m���l�$Z�T�w$9R��8��`���9�~��ၖ�9�$BO��\�F��s4��Ƥ,驧��\7$kW|.kr֌�� U{,p��ބO��$�=���L�>\c� �r|�Wq	����uX�I�~�ƉT����.G�,))o	z�� ���[�³ɮ'aPL�C!<22�I�����~i�%E��F%Ͳ�	��~ˠ�>ݹ�ɐ�B�sǊA�'�1_��l��z4��VYa�Ѳ���uĈ�Tl�~��bS�82̳C��FkXD��������X�����Y����2�^��0j�Vo�p�P8�F�9��5=�S�hg$9"�gf�Q��n[�ߛ[�9��Zc�vx1G��X�B��:�^�,<}�TI����V�bv��]=�b�G��Ka��I>�X�G���?����;��jl1��i��gRx�༖+Ҝq�}7�^ߑ��K �֋6�?�Y�|�~�l��t���_�̘0�Kb�L���+��x�dʖ�j�8%a�T4�葞N���r��BC6�a�:��}�u�p豧KM{��t�3
ǭF̝������^�p�LC���qp��f��Gb�j~��S�Lg�`��H-��c���D��Ə]�{���1�p�c p�ޠ1��R>��`�l��#�\���ص�������c�6��c�TUU�}NP��(�e�F7�C.l��FӇ��`ڈ�F�#;���ڞX�'��a"���*oS�Ǻ4��_�6�T�zJ�e�T�p��I�+l���;�_;�Os����C>B�����wF�&(�0g��2f�z�FI/[�:��u�]`����H�P}Q�^�H����;,@Ow/X����T.�R���@���1�E�qx���|Y���H����Sj/Ez�,����_	P
v�)NA�/Œ�"1�NZ4�KhVt�D1l%ZO9\m)���۫J�����b�P�����0dTD��  0v,|pM|g�۽�t�<�l)��$�&�ܛ?fW6#����W״�5@�k�q-�f���n%�5���f�v22ڬն :��_�U���Iu����J���d���Է�Z�MY[1�jP6�o�	���J�@Y2c�h�Vo��d&N� |��G��@+y��ڄAk��Y�Q�G܂MJK�n\87:	���/X�.i:�XV�����4���*�y������ħ�̟�� ]�k�Y\���Ʉ�^�/g������M�8��Z_� ���4��2�B��LPM���0☀U ����*���n��Q]�M�7�H�6Wt5�-.��<]�ČRS^H��?�J)i6|��4�#=j�"��.�X�������6>sS ��z�ߐ����ꀆ
�Q[4��:����8�|�����`h�_��6nJ/�r�SM�8��v����Q�@N��SE��1�u�t~����'D�ϲ��Jc �F�����Q1MN-U�ww��_�Q��K�Sւ�]bڗ~ֱ���)�͐ۇ��2�W[��Dg^�ԩwi�"�-�J�	�1�(�O�U7b� �5" � ���n��Ԛ��4A"T�l��G���/��z���^����~kVS�p�8���&	���&���]t�iW��b&�QVɚ/���c}�:����&VY��6>y��s�"�8Y氵3��='�t&C	$"�<<c�%��_ܬ,�-�oEC�����8xE$Z1�'��5Ml	���gge4:a�J'ܾ�?��kk"�����f�ޥ�G���S����NI�
T�:�9S�py�4;��x�U���W��c�,r�bۧ�E�>�R���zz�C6x�w[ێ-,��Kd\����n�����M���0ܒbl8$�~hM�͝�R+�u��#̨R&џj�3xy�ݼY��B�ЍcdI&1�@�*��:��Ĕ��j��ֶԸ$��������5�5y���ޗ3��R�z����X\%�'5F��4	��Nt�о�6Bh�'[����#����5��$���-u!#6!�ڱ��|4ݢt9CT��@
�&�*�ESM@A�P�����O�irq�P�KC��<#W�DK(��6>�G�-1gcR�H��vY6�(��N�l����J��
yD+	���*�.��oU�|���f}(]X��a�&-bL�G)���yW�0]�?���o2�����u�F��N��{ם�����ݯ�es�ª������Gӡ/xW(�b;j^�h�c����i��lo�>F��%��]��7�R�n�]�K�է�	�%���1W�<�9�X�.�;@�����yQ�%����t׷�Q��>���(i�ִ�rQ�[�-K�z|��~#H��XI�(j�@�Q�%�\�W��f�M�)���1',�*�W������g��ۥp�D��.q\��o�l7�d�e�>oR8�����Gp ݟ��5'�PHik����[��%H��S�Gl#/7�����ŉ���0�q
b��QH%X;��Nr��R�-��2��l��ʶd�ڮH�����ʙ�D����lW�}���skkkk6�!�'P͛M���b�W����v��Q �7�g�RN;\�s˺�ʧ�e��U�2F��X�$ȿg�8AȨԸ ��!7B��3�7jR�ؤ������nsfT�aכ�q��ԓ5�6 �-��s⻴���#A�	�e�����wE������%�?N����G�S�y�]�VeuFr��wD����t9�eP�i��n	��q<ҽ�d	w�;�sO�u�
�qdh��o+�ړ�G��kOI���5i�n���
�ߘ�h�%��}�������&a܆|�XSN�Ǣ�'��@ 	@-d����L/J�`�b����7w�����_*�g-]��2x���r�K�KȤZ�1g���=-�x������j5&��[C�����3�e�U����v~x����P��3;�lqֆ�)]G"W�ih�a�D=�9{��a�e\9�)���33�ڒ�D�og�U����J�JY���f�����4�mC�l�	�����?X9�J{܉���)�G)��!�k�ٻ��4b��S=� ���������X��_� �]�����P�pyI���{��I�8�,���ϣ*����l>�P8sy�6�
:�(s����e����9N|Jk�y&;���`����_�"�d��U���hfs�+�3��"�Z����L�<k��OhDǤ���b�Gnh�#�W�l;�'����y��1?��n�"ǆW������*��L��G���f�-�Pܶ��J�92r�	��������E�����~S�M�B6�a~����s!7�WO����k�Z=��4���������u�����>���+�����E0��}/�����yі�b�e��~�~fjUˬ��	�u'&���h��_.h%�7���>�/�Z-*���0���]�=��#��z�3Ѻħ�����n��\"3�{:��z�P�<���R�ؠtS)���v)RZ�'����+���N�D�jD����aݡӹAͶ���o�H}`�k�,���=�f|5�כ?��|U�3���ep�fqΟ��>?l�ª�U�����
�2�ґ�!IX�h������3�	�zE���޼�CLZ��VS��H&�=�z;��	k��[-+�DΞ!\��Q8F:r A���">w'���%��;Δ���㛽�T���3��������vJK������ *�0ׇ�c����牡|W�#�Dhʙ���[�[���~E�����H����]�����惟[6������|��I *�X��!}��4f�
VА?}�Ha�a*��V�&e��!����"��e踕KAy�G�B����*A�9�Nl>1@�E(J�|֘1�b:k��DՍ�^7sγ��Rz{�g�~�8��m��9|�>`R>)m�:��g��1s�?�|�����c��z�M�����0�Kob���7v�K�s�_���KQ}�*��vo�^6�t��c���X||�Y�4 ����;2W-���/�j�D�+l-򁅑��i�~h#w��lC��7���ں���J�x���tZm��lZ�x����w�dm�	���̅�מ���?u��y��
6ޤ��e{��"#{<��2������D|���x��(�߶��<���-���E��g����P�*��-�q�<�(���FQU6��.����ksD���;ܰ�ڑ��4��Eκ��mY�|���>��^i����.��[�/S_��g�w=��?}F؏��8�2	,@��2�U��#'��Ӻ�.�l��K��nG~۾2�o�r򔩲Px��Ij]�9:_c
7;aM%)˃�N�	��С	�jY1��j�,a8osj�&g�߷����n�z�pfa���Q#���t����#-��5H�Ԫ����g�Z.��t���7��b�ds|��y�b[O�n����Kvu۝�\t�����2_�NWy5�0(6���(�	�D���js`���>o&�p��lt��~]�p�z%P���6�ۥ;�j�R��O��{$6�����S&��>����u?!�l��V�0����8}�� p��Ah_}/=�P�:ш�3Z*"5�H�
�Kf�u"�IflI��ua]�S�w'
�m�	���g�d$�*�+�8ϗH�X��� �<��}��
�̚$#��IE��d����8]����ȽD��~SJ��k�^�r��!a)(�eڳ ������� �e�	�$���(q����\Ѱ/��vs���ｹv����qޟ����y�3��D���lџ�z(>|.�l.Y��ʥ��������ь��C̖�5I11Ȥ�̡u��yŭ�Ϗ�j��	t�*�j�������bwG*hQcD0���A
��O�h7�5��2F�Rͷ��2���AH]Q�q>�6����4��z�+����5��Rr5��?���i<p��y�RP>�/t$<�|���o��q�,�zq�k�WH퀡6jgGH>�/BwҳD%�R�zeG��Z� x�"u�ދ�#�!�IB�����wg�F������L�ǉ|Xԝ섉�q>��J0��0��Ò��KJ�h>J��=퐾����H��"���`5���#,Ճi����dՔ+3p1��r��k�JM����.�Ki�>��!�7���W%�+zP�4r���S"V9�L�����_r�6��:�KP��=5ɬ��7�0������=	1�KJ�*2M-�r���h�z���VS�cwpX�h���ty� T{_k4��w��f��L�$�;,E��6j�:+�G(]kn����H��S2T׼��s�=p��_�k�	*\�m<��c�2{���{S��Z0��$��ua��D����⹺ay	D�H��0H�h�0e3~���ȉ��]�F���*y�׻�E�ͦ9J����%���-aˑủ]�{�8�I��T'>1}}�����]ǯ�l���5*M��1{@��sVA�=m��mX���g__�?���)I+]��6�q��EQ2�a�0	'ʸq�N��V$5���om�X�n����Z7�{��ʲ�}^���]d����^�׺����J����.ϚXkO�{	���
�"*f^�=܌gҌW]k~��7�ц�S�J�R��9��E-2��a�r%b�����oPc�J��_�"�OM�\+ˣ�g�]��Ӫ��H�7]ii�&Gt%���r�|�c���l��0�|�5�2�ҝ�����wR�2"d�KQ�pZTk�arF�r3���?��Jˁ�.�b;�n�ʈ��	�VBX��!]�/4��s)�;�jsC\	�V�׭�|/�	?�cS��q8���BҮ�[��!�㯏��Ms�%c.��x%!�ӹd}�*'�h�m�0�lBqT�L<m�0���{�`0�{#¬Bc���e)	�r�]����>"�(z��p+|���`Ɂ������:;���`:�&gvTd/��rnO7uu�iN��r�1�Y����{�����jS���A]]V%MA�bA�������=9湞�����m�%�|l�)�o�2�v6F��]u̳�Z��q�#=� ��L�,Uڥ"�謅�Ň��9Y��;p�9H��_l�8�����ǐ�9<��2���I�4Q�����;�L]�j�Rz�y*�?C.�/���~V��a_������/Ty!�ѶA�k������[�������D'�s�آ8NICz�.�o�#�0Q��A<�l�٭�ǽ�{ާBgȒiB���6�&���ô��w$n�`{7���Y��H0Md)%����u��O�Y�&�	ʶ$N诨L�xu��[�����nxǲVt�Un1���YSn;6~-t�І�{>�
"��ݦ�Ǫ��Y��˔Y٘�>K��6�iQ��.�𽼍� ��V�5�W�'��[����� �˞dN�b�*�+��J�v>^	���]亸� �����fG'ǒ�]�*t$H�D��
�w�1�&3r/Js���-��]E�h�Kk�cX-Տ��G@��(��fQ��:��Rt݁i��;���5�?�\�`-�,yˎ+�ȓJrYmi������{�v<�����_�ToR���(	��>+EM�dQ���DN]<:T�B-D/���]�f�&��~ZS��V��)�~���a.�2dhnQ�O�)�N�9�b��d��Uh��;:��B��m�d^�`�\���ƄF)O�0�pu�mU+���Q�)���z�Õ��'�|��n�@���]Πo.��'��-`�
3�����v�����*�Q����������_9lkc4�����7�H�w��q������L��Z���1k��	rX'ujQm*�����p�ԗv�n�HK�N���$� xĸ�׏biHL��R�,��{©>�C}6 j�.�CRO��i���S�[�^u2�T���*�]>��2��v�Ē*7Mnh��罴�<��0��!�eN�43��q��s|w���և�<aU;:+gZ|�l�.�-^M=�h���������!C����d�,�n���%oL�aˤ�V��SЈ����\A��A[�=#;S�V*��u)j�d{&������C�Ӱ@��X�񌂯���4�x} �ҘP�:�<R��q��^KRW7��l��`����Ѯ'�<�?�#��lˋ7��#�l8Ց�N�M1��������mnv��pv->�#x$�6�-�����M�c���v�2�/�����s�$CƑ��&��vqjT#���H�蜃�>G�YX�9�>���I���0c�;"K�l�U�3wj���.&�g��(~b<6HJ���y��SWI)
��y�J�n[�*��HE|�Y���}�����a�:��7��c8��0���Gɤ>Mq
���=L�3fH�A,�_{.)���O�U2TX,�Q+4�L{��+�-<�a�Bo�4���iy`�T �^�|�|��dr����j��0y�\%�@�l���nɭHP�ds��=�*������qRTd��2kS���6�h��%�t@��[c�_�A�D�\�,wX��=4����V��� �(���&,-�ˊ�c�+�T��,cX���~hO*�\�:v�'O*>JҎ���x񮱃�sW&��1�R��·���f��wkB&�%���5�:t��:��ZJGJ�юS�
�un�:�����R��i�ҦX����F�S(���[��O_�Q�>���3(>G���(���YSr�	?�
� �EI���ӵ���ܲ���`q�Q	�T��XX�X$ ��O�P��O�7hT�i�D��\0E�]P� ��F$͆�v�KkB	:[�*jKHPM����Y�_Cr��.�+�RF�D����f�dxNO��L2�7^�L��.��R��6��Ϯ7���X@k��i}��# ����u�ϕ�P���h1��R�^��-��'�	;p�qL�+ÌI4l7s󦃭�jl�]�kwY��|'��""�L8k����-�F��FVi�-5��GUH��#��C��I�*�/�st6%�KŐ���*�����aI���Rg���[%�p9�řx�=�;����=@��2j���ǅT��/� ����)r�MD%wi����>�d� ���(±8�*�k�X9�IC��
�X�/@G'�G���j��sA�Ż$�x���KkJX_�da�|�YF�:#[~�j�LU������'�-E��6�T:}��:�lfU�.UW��<���	�|eڑP5:�o���Z{s���TTA�Wmqi�O\nY1+���U������V�4�ni�;n=|t��E8ʊ�u�U(���g���D=~�p�n\Q�8Q����#�A�摾!�O���)ܽ'�0o��}Q�Kf#(;s)�޽¢%����!`��Ƞy�Ƨs�W		\
��I�jq>�;H�j��?R_[��,	6vϋ�Q���z��0���1ש�O�Xb�'�4�EB��rJc�NH?D�2�Y�Vm5���2)�6������` |Х5#����rC�%��X����f��X�##s�Q`èqc�,r�O�Y�=η/]vC�e��ܔ��Z�z��eJ�6e��P6z�(���Hu� ���ͮwK�k��r���087�������c�l��M;���-T�,��4�k\`O��+���>�.�ub���Af%9O�M|6[��Fqxf7)���8L��@��+�yB5��As;m����<��N�3�Ye~�:=>���)���)��,Րէ�(���Ώ-"����@�G�+T��, �
@t��9`��ذ��|L%�\�a�<��Yo���UW����O��]��Z|V����Wu3b%hg��eЃ�M���Ν
2��m���s6��uq�qph�&�Z�i>|z�EY��j��N8S�瞑{:���b!D�9}�xLxUT�pR�#\6+B�����Ӗ�R(p����{�`���d��^��tTAű������*�Kz��k���즸QG��˚��	�w�I�jK_�M�	���M]�
h<�_>�����I�7�k�{�����a��7q��5����D=���]C$X{"��Ko���"����J�%ޭ��O����-S��7��]8�ċRv�`U%ze�\�|*a�@�b]����h�"�U�Bv�HHF�����m�@��:�4
�H������V��{{����,O���1�=7Dn&�C��M����N��T�[ݼ<��o�xf\�E���nC[vUW�<Z�o�$(Y�Y5BzT���&�,8Bf� iq҇\dV|����T�6f�.I!�vf@H�i���"�0�x@wg��4�����Cù{o��9(P�e����()d��2_�b��Q�ʵ.�6�a��^?q6k43*\@�i�D<��b� �h�ڝ�gX4�䡿�^E��2��kf�\�?�(�xl#Nuy����5��eJ�&� 9�|x+��tH/Љ/*Z�^aTy�}3��o�<V���d���\8{���?��o����� �I�3a^�a�4�C������X*��<E���A����!m�����~DuoL(cC�)�6��\(#�@݃jDW��#q�e�ke��D�d�g,��᱕~U�� �����J�p�rF���h�\�F��`��f/G�*Ɏ����.2���p_ﶃz[6��� *o"���XN�^������*�9�����q�yϻ,�
3o�>��:Pd�d/yDڣ`3�ց��
�CV�]���v��uKm���
f����iږ9�9y�rt�������Q���o��2�cB��lH)���|�KN-��j��!?�N�h�ؑX�z��%���	�o�J>���?�T#��������teq���Ɵ-��fs���$6?���#�+ 2��=�ne�W�F���x��Ƙ�6	�@�B�cX��� 1����耆Ɩ/;��2A��]W�ι�B����+D��ؘ`I����]�m-_v6��J�����ķ�E�	N�?p�z�N��E�E"�~ݢ=���p�����f��U�J��1����.��=Y��G�������ZqXeL�j�:�X3Ʈ�/+H%
w��PAi���ތ�#qu�o�Ez�t4TF 
̃�+߸�	5G�m#�1����ʼ�m�ѧ�����z�ԙ�FKX5��(��C hhӽ\�Z��O+��>�_5������:T�l܄K��G��t2�Tn���_�g� �b��`�|Q�'��������Ǹ�0D�%�$����1�6��N�:`���r�	����-�IL�Z��9�o� ���~���
��{�/�T桶%�ib�S&1nIt�p��v��]_`)dΐ�R���Ŋ�U��;tf�[2f2�AgNc��ʬa�iL��y���{|hR���=x�I1X�o�n��_T�J�͡��CE�|�{�>�E� �<��KH��D�o�G�	D3'ѯ�5SA��[Bz[S"}^�m�ݮM����T {,�`;�i�o�Sg@a���ԕu1:���҉i�Ǜ��nGL����P���[��O��X��<����ݲ8����C�K���#�'Ƨ'����W�Ҙ�Q�4dX����[Ԉ`�5ˈ?J�im�[��r�;wmHH�[��'#�HLř�.�9���p�(��@?S���׶}���O%$I8�u.-H]H�KQ�L��-����}������#_?�տkU��CI��|�"��%5�) )S�f���}�d�@�Whh��>�z�����ɻ̙}� v�g�'w����0�3J�%U{� �O�D�b�sߚv��: �ö�j��{�Nhr*�*M$0�G�-��3}�|��s��4�
Y�Ԭ�A#��I�bc��p�5d�零�U�>�CIm��t�3����g�Q�솏��CLt��@��Ғt�9��&@����{@��ʱ����v�^��)��mu)}�O�0���+ɷ�(�i��ġg|�
 �q��n��'4
� �����\�]��y��^�޲wM�!��� B�X��8ڇ+��i�eő���;cgS7����-���L5��Ѥ�٥ESS��,�l�p�}o �ӟ����E�!�h	Y�vn ��
�&�[�G!��+��։�czJ�#��Qm�0�X*�iٹ+�K���i_R�^:���V���*��B�����"��:�
0u�lauy�c3g��VQF0a�Y��k����3{s(���\<`��s�Hq�����!��A�}!���_�1@�}�C�]�;o}a�m�܋驴�����k��M�=7�j竑J��+��&��E�v�Wl�ݹPu��(}����
z�*�[����L+ە��2|�m�al0?>B�1����o��(�Ud9��)s)�$@Mq�����13{`Ĥ���]PY��0b%��Q*p���#M�*�I"�Q�?�K���}o�Kԡ���'_��n�~�Ź(�\1�9k��H�H��l5��U��*tQr:�rM���ĿD��`XBBa�C�>{p8$�6 �c|���U��_�%�֓��	f�K�׊F{���7Z�l��w]���&i�ضm''�m�67��ضm�Ol����qǸ?�a��3��{�\�f�iY����L�&��OP�O(Ѫ���39�I�,Y��)� TCՊ�0n\n����|�G��<�{uJM�|��!}��'��f罌���?�t2�u�U��%�L�W7��V!�L�,�$�ǬO:��y�q��r��uPY�<6���e3}��F��$���w�'l��LD������R�Yq��]���Bܱ��
��	��=>���X�M��5* @��qX�9�5)��3��%E!">O�����_0�7�Y�_�O�P�޻9V�%�(�������M�k0�%'$M^nv^se��>+�%�,q�����Ǥ�A{��҄��D�V�])�%��ȏ�-R䘛�h������?Ut%��c��6�S���	����M;�إ�$�D����<�Т�k`�D�X�HJ�;�ֳ�$�XE��T˖_���6T-4���!?11�2Z�7|�Y)�k��=�&FSu�P]���*����!t�������U�!iaS��
lX��L�Tb~E�@ǫ̓��3o���Q�K8�������	�~@�ߑ�PIM`5�g�)��[�w�پy��9���r�"W,z�����\��ݚ��|˹jlh�v�Kkq����CVY���:d؊��cu�޳���˭W�n�ohP�q�٩f�+�)nk͞2�8n�݌^���O�SHD�����}foaR�۾�{V�K��?A*��6��D��٢r\.����	@�Ǯ��+��T��0jQ��i��%vP��L�hgmi�rZ����qG�FZF^�yn:I�60�?�"�bAH��Y�?���-$���
,`��>����_�U�._��QiRQ�d%
�r��${��e�٬첥���ORTA��Z(�6�&���`Äz�>#�ֹA}h.�H��u��ޕ�2�9�~�.�!y��g��V�>|D5;e~~<o�ٚ��K#��n�8���-Ϡ��$��{}}=�?�'QW�����tւM ��L��z1��g$[�@5~�)� ����=��pbCbX��'HZ�\t>)���ot�DGˎpĚm�ʙ�0�-��Wm�F����5j>���K=1[�z
p����)	�"]\Top�$�R���h䪡^�F���'���)��v�:��Xuo�À�E���d��m�䏌b��#�����b�FP���6��|���$jȊ����-u��'E�;�������K���1Q��J���<5q�-bǑ[I-Fs1q@]�I�ȩ$��@=b|��"��\�C�#)#ݚVT؈zw`������ew�k"JK�`��lEIMWx:����62R�ͧ���i�d�x�5�~Ӷs���� �AG�szz�9��E_�;����&LX����,���P��A|��$`վ����y�-�N�Ӵ��*h���m�+u6��l����ڬ�C��$�R%D信�Q�>Sȯ�B�U�%g\������u�޼"v����l2h�a5����&�����k&`AE�%Ct���ڲ����c~
Ȋ@?\����⬙Zi�ڧ�ן�QB{*S����?��}O��%�G���߈j�.Pw�=����k+���=>>�����8��$����M���+/D�(s�8��s�� F���.G����ȕ�R?]h�N~�OY���2�{��(X�5$�c�@��[����|���9Mb`ɩ&��nOHСUU �(AB�������e�ln�����������4e���+�촱)�^;d�qWx0�Ijv���#s�l��qGG"�h�`89%��T��w{3t������j���=�סl���P�צ7ϣ��{�R�sI-X~�@�4	o�e�c�wgѮ�#i@F1TB2�fz����\X��/�V������-�m�hP�����ON$��es���'��0�\os�j��B�.��Ǘ���=�����;τ�jl�EM����B𡙑�d���	�P�`���X��|C���i��i凤w�|��y�
"��8�$L-`�tb�����<����͟����\�yWR�l��16���z{�*�K� ��/���
9�����3b�4w����Y�{*wg����o�o
G�Teܵ�߶�~�7����w^u�x�3�Rp�8��6�ә���-�	-����Tc��p$��r(+&��)j5:�s�x��M�󺏟���Pp��	Z�0;/����W�]�WK�[��I���AВc��W�|r5z�$e8�7v�r�l����"��Gi=\�V���Q!]T����� }�K��>�ӂ�'�NQ �߾��k��E���G�����������b��m�HB�����-�*"ת��/�x\Bw�S�%I��xӖ���hK�"���6'�ʗ��k��C��A�)��!�(A���.�R�`�)�,O��8R�I(��=^�_�BT���K>MV]�<T�C���� ��9��!99�;6*Q�����
Q��-�������W�=�t��8͔�q�<�f�/�V(Қ]՜"sSeu��Lv�b�HHؼ�ngj�.E��Y~i�ӭ��9�F����.�n���e-��#ް��	�"��s�њ&'�z������>�+����X��j��|�@0){J�̑�F�y���p̨���k��A��HU�]!6N�'"��Rؿ�y���"N�r�?MW�:��[��턗��]�v���Mۏ+6�l�2��Y�"��2]��HqM.>.]Q��69:����)4Ƅ��u��G&4ҥ
�yLxo݆vj�8���)[{7�����AG�{�H!{u�T����aH��rw�n�W
��B|�bR$��2�u���
�e�0����PQ�5�/AQ�S3v÷�ʯ�ƚ�@u:�z�z����"W�����r�g��KCv��2��Yb~s�nw��9II6cw^Td6�7��cOTF�Ĝ�^��25?�r��cqZ��ȱ�km�M?�o�Bm���P���1�_dJ�;�8o(%s���r����Z�S p�I���&�%��;�n0�KD��H;S�
;o(�^YQw]Ю{?� �|;�i`�?kw���������|ʐ�9�H��^�D+ƣ�F�(��u�#�ܳ��������r������cE�
�7V�پ�YR����t�R�j+��[dgsl,N�Zqg�-Ȥ�8[���v��S���n�~͑��됼�j��ǜ�gB�y|C��Gn<�~p�|��Z�-����PP@���x����,�{�ٓY!	�=T�vF5I[R��/���g�N�=�6���C��م��5YL&M9Ig�)��V�'�` �w��l�X� ��ue�\���*ܴ�g�u�X��veU�+��,M2Do�5�joT؆7*���@O(�;�	0�Ȑ�~מ��A���0\E�7>��ŝNo
�5�g���R̂������01M}H*)�U|>�2���7)��������_�����i��Ƞ���Bd4||q֟�+���qkm���N�������������A���g]&w%;b���M&��Z=پ7���l�p�:��͋�~�	���?hg�"\���X��Qojq��������8�~�����%WU�3׌��_���~!H�\T� Иɣ���� 63Ƈ���M�. ihh�p���'5X~���D�h���؁r��h��\����<�Y���Ҷ|s��Sd	X2[5l�89���F��
E�!�>�{tN���J��'���;8/��p]�Q�o�� ��p;V��<#+���1����G��;>d	�nD�
Ew]Ѐ�C�K;�Sg=���lH�;��!�������������B�?����������N��IZ����n��O�����O	Ͳg�Gm�#�\^��}�IQ(�F�����:NF)Lӟ''#��������a!�28���,0�w���Y؃Eu0�s�8ѱS$�qV��>�!�ܦ^gV��'���<�9��9�����\C_�� �=8� ��*���'���6�_���g����k� Zi���P�"�@��r
mkGAI��Օ�uq��Q�հ���$�W�w5���I%u�7�Α�ey,�b2J;R	6��99R��o�Xj��ϯ	��Sٺa
�}��P8��� ��wB�)��:P��BL�i>��D�K)6GC`e^6��FϽ�4d�M��G*����}��H� �$r�h�10�����z��1����!z*ڶI4��N��s�R!�״}S��Ӕ���*]���&I�I��8���'
s����9����]	��<�)�=NeU+���YvSasb@�b��Ǭ�>��w��e����}ʲ�d|�@��6�OOƭd�cH\B�B�<���S���5�r��6x�y�3�C R	+,���*]�-U�lݭ��\/H��Ư6l�b�B�O�G����灨��n�}�`H��_�mίl^��U��-��+� ��b�'Օ���?B�����Sd?����e��&�M��� �?]u��-A�����]��XJ��Ea�UZ�������iV'Ǉ��_e��w��'�Z����?V@�OC�;n���P����4��h�;��%�^q�_ɖp��H*&��9?A�}�	���#�v�\><Z�^M��;��1�7�;�ĮW1�	(�k䭌������S�]�Ŷ��_�;ۓ8�5D���<�M�n���T2�U���/ONR
he�4E9-�w���K�NL���h$|�|��U(����l~��D�b��6����0��<�{gf=���i�u�8���}l�9��z���_{P���8��|���Jn
�)a ��R����8���w�+:=q����@D�Z��+'��!��Fj<���`�r]31lܴ-����B/���쳞+[͎��ّ-@�w��=�S�#���2<����&��Q�;	g����D�>�L@�#UP�H����
�e����5g
D�C��o������VD�=��h�a��]_�xx�}',��ʍv�g`��$�0��|�*���vx�� v���Q��VV��p��}��n���6:��#	e\���6�J:��8~W��o��$�H�%���}����cT��惕Sc�6�����՘�D���[-t!�/�'�]�L�<��X\��&Zv,D�*�gщM��+�μ�٪��~�P���\�4z��{? ��G�<�s�W�Ŭ� �^�DhG1�
��q|�>�5�mm�+���s\o���_`[����r�;�ʺ���nf�ߗ��ngx��W���ށg"�WYw[�]*��[��X<�	/Q�W� %x+�@�0�`7E� ��(Y�բqw�k_QIcr������
kJXH����|�TC�;]���wSu�XS^VT]S�J�+�|��U����ݝ�Q�*���I�9($٦���Ab����7�����G[��:3P��N� =5f�q�I�d�n���=Sz��
�|b�X�Wk�]���s��뿡� ���;����X��P���+^i��偑������Ğ��3���$J���jd�f���{�X���c	��y�e��"��Rk� #���ޭs�s�MF�E��e�B��M��i�W�� �H�b�,�T��}+�m;;z- 9�x�~��\�����B�L4�����gɴ�~UR��$r��Γ�����q���:4uª��G�2�i���5BK%3 �6�E�3�H�Mt&HwTn�+ثS��gs{~>2����x�ZȳZ�{v�$=q�[�2��M�C9��= QNGA�DE˿���\78)�� ���8�X����no�쭈	�ƾ�~	�������E�*�p  ���a�_\�sX-b�n��(���Y���H�o�i��8�����ˊ�`#�Z}-/O����W`Ȍ��9�D�|n�8t�,h�::�o�낄��l�(8��rY�IZz�����
�N�{���Ŕ£/2�n-&8b�6�s����Bp5�G�w<�h�윬�X�<�\w b�K,��C���2�B*�(�� �#�ɳ������B�UG��g	ZZl'�;��t��Z��u��$��E�5�ݙx��@��r������F���x���v�:�O�w+j��[��p�A3�م�
Lֺ��z{s�zlp�!���[IF�dfe�LA�\�'^��h��,r�IC�<	����!Wn��;�>�����N`ӃƬ����U�C"�a����$�P/q�|������w��j����P����d�"�$.�����>�t�䂧��*���g�]a�`?n�"�RSs�S���ɡ`bX�	rD��~Ub_���5��	�n�X
5��� ���<V(���j&�v��o.�dĚ$�x��-CC1ry`?ho���������|QMCECe�{eYMMo��e��_��Z�~��ggX<]�b��J��0��^�o�^�S��Qr��R��sV{Z���Z��p7m]�0��J��\g�6�ۺ`�i��J޼Y%b�������b�~��~��c��l����Y�+��� �F���%W���@>��hE�b��0�Aa1�1�!B�b"�x�ƧaM�M!�|��5HZ��(N	�W0E����?�{���y��,�N�=���{�[����=r1��^B��HD��&�_�[�;soo0�P�
r���|^]�Z+l|��`������D������s�$DoK ��r���2��P�
�(���'#T�����gT�)��_�����&6��-o�Z��H��2|M+��-)'-���h�W�E�
3�A*��O3H8��1��.� t1r�,��Z�xU�P��	��3
�%)6��=�?`z�+3�V�To�Z���c��H���2�o��-?69�D��M����K	�
a?WH���w2c�Ԕ�b�!iݮ""��]���Q3�7��O�d9ݧR�(_��$��m��1�$�1"��m�vS��a�T��T�!�ϣ�����Z���=�'�F]�kn]��RV�q\O�j�
�i�r�o@�h��|��JeOS�+����_94O�m[$5�W�=���(�B7�ϸ�$	Nd|n����8b���U;o�opy���ӫ#�]�>�~~~pA=��+e8L��+�g��քݜ���b+��Q��l�S5����mQ�U�/����	9����!mm0���"�(�s���)�$"i�͚|m�;\�@�Y��4�i�e_���;utSDq�Ʈ��]`{�zA뺘�?�z@|���S#y�+���|����c�n=�l݈y��S��6p�d(1 ��U�D<=V%TXiM!th1�H��6|���+�*1q��=2')�Bm�8�Z鹒$E6
�霓���'�w~)�Ө�����m���7\|g�4�����d�X��F���Q�U,%h��5��]��V��}	*��7MP4[C{�DiC�0G���@Q7Y�F�����Rl�m	�#�W{4��͠�����QȠ�<�[�m���ݏ�罸�Y���v6Jz�J]��RĊ�kp'fس���L��"�4Y�*�����v1,��=�}��+"e2��#��V}j��uF�f�OH��鞺.�S4g���
H��i�*�v�=oV����Jt%���F܃��gT��yLj�����J��"Ԍ~�$0�� h5x���X ��?��ڿo�b3LL5*
��Pn4�"��Iϋ%����Q��h�{
���#7�k�n�>�Ǖ��_}�t����x
�A~�@�\_[��#(gվU�py&�&���!mod/���MZ�a88Rs1��u�>G:؊s���8d�ZB�r��a<�X >b�����D�����.Y��r����5�|6+o�{�j�/��"'���@h�:��%��Fy/U^k)K��2�y4��~G���Nu�VbjB�����g�6�KV�ݰMyz�;E�#)E��E*}>C�g�4o�ލ5�ؠ����mC����~Q}���X�D]g֧!"�.Zj
���	�Ě����w`r�a|]Z�2�
���tB&Tں[n��;���6Ҭ�6hܦPSɫ�ҹ�F���.v��������A;�������w���{8�)���cZ�:��&]͌<qA�f�Fp"CI�lP����ƺ��0��dA0�:N$���격2�ԧ���(rɊ[�H��7yx0�ڂ#���$�)gkz��#���3f���5��8 ���(�H�zfY"?�����T��ɑ��p���~��Ϝh�����&��5�����zѓa�U�}�(\���Z��j+B���ʭr�a�sZ�o*hry^ǻ��(��7ip˥n3� �D��8A=H�l�,,'�6�h���b��%�CkV�$��$8�Q+�{TԔ�x�+7��B,}̜~$#���]J��2�C���S6r���yK�m+$8H3��*�!�����3��m���˸��$���#���ٶr���Yx��M������1N�}ĝ��.�=Zޔv�q�(X����B)���o�|]-�N�>9�/�W������Pt�(�����ыZ�9�Հ��|�Ҽ��|�J?)�T?���Q_ �isYI����y���	ڀ�-�N"a�������Yo��5;|׾���?#X��s{������Of.=�4����z\�7*�����$���e̥)4���s�D��&{�xǥd$��#��Xm*к����V6���h`�xy��/#���Bs�	�0�m��Ef��u }��-���Fe��8;��9�"����;�π�]�
5�i��;�"9���cad��?X�V�L9�93�_��!�����}��c�SBn{>���N0!}4$ !����Ӳ��/���ëq2��[@9�颏[y��
�	G����vYv$逘�걊��7ctX��MK@��f"*���c	�'��1 ���Bb�����Z����?'PZ����iT,d��?S����7��FBe������q�%X��V�,1�_�����9,�Q��R&�kF��� R�T�Z�-K6����F*=on�S?��a�2���f�(�.����|�D�;�Y���!ASb��_ۀ7�q��g���$�wO��j�C��"�B���q�B��b��ם����ωG��>�	t�c�[&�ef�Z���
�����'>5`��YP.�n	-��^��Lg.����,nI�sbΒ�I�>�
һF��q������x�O{�n��B�j�|��qy>��k�$�:�%Rdh�9�B-���2QT��2�0ޘ�-&N��J��מ�ݹD�7D����}��;!&���"���FGO��O�6]GXV�����Ke��C���J:�I�~@�@E4���ۙw�l��Qj����ѷ��YÓ���W�V*�m����/�x���:-�{l����Q�a�;�����捧ɀ��K�0�h�lAQ��Ć��6�>�s9|Y�~c ��h�i|�붝�Pg�G&�-"�a8S�5��+�e��+�Zg٩���������㠱kI`3���4ʐKx�
���Z�C��C�����)�P�l�,���+���l���|��ѭ�����9����$��k�}�[�k&N��>"�	�L�tx>�uH��ߕI���K/�Yn��zpi��g�T ��"��Ο2���
>D�䝩s��b;��G�d���(_D�X(������#-�w��f��*_�o/����8�,��acP�7��*%-�Lh�6��p�W�_��p�rr�{����Eʻ�%�
9�}�S�7�-K��n�95�i>m�4ⶏ��b�l��uik��#&����:�|����GyلF#�䲿�t�K�,V�����ί�f���k�G�����L��`0\�0�q�#���g��:����jT҅�e"�G�eK��b�c���sa�N SA��l����Ŏ#�`��M\c�(���n
h�t����ڇ��]��i	kk1g��gh!���<����2�6�e�k9�������H�o��{L������d����O���_���<O�3S�q����NF�!
�������|m=�qI�eB�M�X�c��Ǚ��~��ͯ�A��.�LRVp��a�bx�������<�gțG��i����~U����4��`�.x�+)�fԀo����:b4�.�!p]�y =�\[����z���21�ff1�e�ࠩ�-N#�����=TL6�0� �� �@���bso�GJo�1|Vd~�z��
��1�=�N����l����+�������D%%���m���L}zY��6
�J���Sb�,G�p4�G�����	�\�Ǵw ���۸U��+�/��B�h�g<q�O�m�{�&�5����O-cT�'��<�Q^��4Y�~66UErkCCfT8��Y��55����3��f4E<�����rg��w.�L�?(H��%��\��`RZ�i�����1P�k7�'9V,i~����n��:Ԏ�t����V�|:S�*Fǲ:�|�������7��`#4ज-��0 ������#��&��;���w�p�Z�,��b��ܖq�����s�3���*!<�� ����݌�OZ�Q�`��c��v�Ȫ'k���B�a�G��p �-�%��<2H�W�C�6;Y osK*G���	?xV��T�L�$�<��1����9{~��5ZlzK���L�Q��D�������
��g��a�3���g�סU/���B�s�E������A�G���{�(��V��*O�TU���*m��A ��g4#5$CN�'�C�O���bec5b�y��Z��x�L���O��$����=!�>P���Ix�����&�go���t}�x�JhY0t#ޣh�F ���d)/��,{��d��g����qs��̭94�<���g�ۭ�kEM�X@��29ex��+2\���8��~���{���tT8� :>' �Y)���!�xl��)�p��pYp�����eh�>.���.�<�;5�Fl�0M���%�Hd&HGeMS����Y_��>;����N�׌�[f�Fn��>aD��
��-�D�RU�Z�|�>ߒk"G��B���ER�?^}*yKJ�ȕ��/�v��$�*b-�h�M����l��+�t��|=_m_�9���!;�M�z�ߧ7$m���G	�4��)����)���8�IQ7�s�QcN�@N�逵o�q��	b*�7�C����(�q��txa��WP�������܈���͌?�O��ޔ���'��x�9�n�?kv�$I�����)d��E���~�"�`��#��&�/�՜�(����_�n"�ĳ�O.��h,�dfĩ}�uz+}.K��o������6��,(y3�FVaRZ�Y��+Ӊ![͖ԩh��8��˧����m��z�'�.B	�)�w�k`q\����ym�����F���Q"S1��(ۊz1GLj���+�ɾƠs�,��jU��h�0͟s��=6f��説�)ܵm������Q��eE�V�o<U6��g)���a���Y���Gr�l��9^)zSu��.�H�oumFѪ^A���n�>9���S���LF,ä5���/zb�{�Ү��������%=�ہȚ���t��Eo�ҩ��L�O�Z�i������s::����Q6��<��G$Is:�-���Q��:#S��̴�z�Q'249�+�UQ'qx�A�.y�����)[
�C_�p�5���7����l�|��s��$�.��P�������}Z�
�������	���Vg�7���93G�F��^?��F�7�Y�ݝRB !<k�3�J�~ak��0<vpW�����Ѓ��=
r�nx�{[^� !!)��l�����n�uѳ�����������$����Nn�S�v��)�Aw4�KT<��X�y�e�+5p�T3��d4L,�y3��UE�Z �Ȃ3�z���K�
�u�Nr^��{r�FW�����899��W��6H��͍�������
VP���,JbFy	Y�>"B�C�Wʱ� 1�mU��xz|�Bf���;!�@@�zڛ����P`�v/E��"!_Sh�`{f3�uoj�g��g?F�ѻ:Ϸ������?Cp��Kg6#��`N:4�H����\Z��`�8��L̽L՛����`g���4(@����z�u������M��i-x�����g!����o�Z����nt���A��9�H����;<��I�6Gպd,PBm�?�[���K^O�����Q��Ⲫ��ҿ��[6�F��nB) jd=r|���QE��χa<	%Q c6�j��,	��֤j� �>+�̶�䪖 `�e��1��L�e�v���v\FPP1+��G���ȿP���O�D���_�&�Y��}w�'2t��޾*�D.���hԝ��bջ'��_?�3��2<���6>3,�NK�HCi#�)L�1���/��u-�i�¤���de�z8�`��3�T_npY����f�	��PLN��OZ�3����f���p�t<�I�69ˬ�ʑ?����ܔ/�;Q�`�$ʦ�ీ�t���Lþ�::��(��'�Y��q���@�`����JI8-��*e�.�ˢ�o�;��]o�a O��u�����gD&G8�ݐ�k�!�����=�3�Y�2(x�AL2�D���D�]UN�F%�y|���:�P1�`!2H2���z�n����/�*5�R��Y)_	%%]k��3�����^� �޼�>L��;����_�Q�G)�9��:b��iL&��u~�ƙL�q&b�����rSD%MO���>�b�e�<g}�5�"*G��L�w��Ó0F��a�`�6J��q|�_D��)�팓��n_�\�=�ʍ��]���ԴT����-�[���8�=�\�i}�S�\)v��&g4�
;�����\�ci�]��CX�^�W딡�{3��6P�����/��qP�Œ,�2�в#���2b��T�a���&yy%i���&keB퀖<�p\��܈����v�]�ϲ�YG5Q���9�)tr%o�k�y��ATS�Ay� }2(-�Ǒ*����T�NFw���}l�u����&(��z�^ӯ��m�i��,`_��c�_�C�fr2>ol+�E��X�.�0��&�"Q��G�vt��D�~��P A�����P�	p7X�]�P�s��/�l �����y�L椈�4�D,aa�Q�Do���V���)�5���`tĔN��7�l&[���rbf�x%��|P���ۭ�:�5�� ����27��$��e򔅽�G�-lPwf��J���6��@?@����ȗ��@�Q@O��8:�ǣNI���`#���`-��l{�x��>�������L�o�����r��))�$�n78�ֆ�0�"bMiJ��RB�أVi[��O�+b3#�mQVW+�������
 �qk]u���@%Y���4��y�'��#�۰���S������b���%V���v��RSAt_� b�Z*Y�Q/P`�D^��m���I�L	r�8LQ�ɨ2�kQ�	G�'�~��K8ݏ���r�d��ۛ���ť�6��Mq?����U�ͱ����39#:wG�EmAN"�u��ҷ2Q�C�U�����!�:��.>Hvh�
��	[�.���˃�Fs�{ÕbY���NK{�b�9�]tڌ^�����p��FIp�A�T�JWJA1NS�w����%��}̻����4⇀�6�h���v�{�ֻ봞�ңٛq���kXK�1ɱR��P�t����se�L�c�|3݌-r����1�h���}�>��� ������"���/JU��2��U'�����?��æ�9����z�ʲ��bߐ(l��:���0Y����fT���F7���J��4��<oV�$��.��	"V|�d�$u��'h���T���=��UZP��-�v�.�6�vD.}���AYUox5CE�Ǘ� �]�;,�3I-}vu��i��>�zT�>,�uI�b��g����q=h�߼�}ȿ0��]J�akmajsG��L�Q:#�VેDB�\y�|q��RL�3���������-L�����s@���j�%�=�����z0��qAL��	A'E�NTn穭x�kx�)W"f�TVlj�
3L
-��>�aLYӄ�L�������K��N?���=Ĳ(Z��� >�}�������т���O��j{���Mh�$V�d�d�������>'b�`W�ʢ՟D���X���C�e�XN������	t�̇$,b�
4�B��P�O}�_Y-27���{���L��X[�=!��S���/?�'�B"�t���0���u87dr�Bc*�A�X|�������˶�=��3��r�%N���<�z&��'1��/k'VX���1:S��kV��R^](N��m	�g�3Ȉaq�o"%�7��%��!��S���J�DM��uz[r{���Z^]JkО��'��.�46���'�1�
`�CdHq��YOjW`p:�X�RЀ�����:�_�t��d"k�(Qڷ�מ��m/�=�IOGD7[/�T��D`g#
\��N.mB�J��X����S%�sr�'Eu=�A�BM��>�l�\�]�QtiI���|�@&��-G���Cg���,*�Hk��fW�����e�іV�)F�՝��g����[2�9R�4I��c�J����������;~��#h.E�=�~�p|lvx|c�Ӣk��L�|��U�|,m����B-�t��EϜ�7�(�߰u8X\S)*~��āE��G����{ζ_x/oj��OM��ۜY������y&)ĥ��QQ�����G��邻e�p��`ix���3�-ܶ�1���[�ۤ��I0"53�9�f��$ ��x)��C05"�`�Q�a���ԙle3x3�`E�^�ډ����=���2�@�S�i�ˏg?)����U�4QÛ��b�cD�x�h�a�Y�!ٲ�o#s��ms�B2
�o[�"�{��ޯ�@��O"o��I��Ӣp����7���?]=2��������l��tΡ�<={nh�p���y����N��$���E���5 ���8Ƽ��Q�י��  =�{��b���W	�s��C#n�M����S�y`n�I���M�5l�ɖ��t��;7y<����|�gD�/�� ���G��74��n��6�k��Y���5��r%������\�^�/�79i���V
�y��ϙ�ΖW���_}���.��g�q��K}~�}�(s5x������T2��1���?�UBםǂAE3*�?�ON��<\8sIXC�I8��3�u�鴈X z��'?2��sao�%���"3�X2�2���?vkx����\��me�����%��<�v<ޕJ��"#����B]���{�l[����K.��ߕI$2/����60��s��k	f�Y给��{vRz-�� u?�p��$'�!��Yt{!�7�oi���Aħ�ϕZ�Wh[��f��O���Ѕ�b�λ���i�KSde�U뽱�zNG.�Ȓk`(����O6�=ٍf��ӥ�q<1Ğ�Ag$~J\ȸ���׿g���l=KǍ�������B�cɤD�!q�,/lL��"V �/��[�Mɐ���@#)AHS+�8�Ne$)�]~nu�,i\=��(��r��8[y��nY�w/럽�5D�s4/e��!��Y���(�9��=bw+��r7zz�d6w�2�@P��w/Ԅyy[~��$�)�^�	����1=��02��T�P�;]P��i�	�Xȓ$r�3b��ҭ=T��}��}[,x7q!��7ԮЇz��6��؅(SX���VN�|7<�?N��<���u���m�^���b�����o+C,�_�Eh�*�JR���ȩ�?r��rU��"=�h�a��Y�D#��z<�r���F�����k�E��J�2�E�k�G�l��H{Vo�]� �`@F]H�}_�{?.�R�~��ތ�ly}���~�d �f�B�Ĥ�}Mq^�U�T%<ϡc�[?��IOᑎ���u��E���-l��5�̱c�t�w����m�OIt��9�SP��3�<PLD�m�HK���j�R��z���b�oyM�]�ۿ퉜s�&?Tr:�-H�ۨ�uFϾ<�N�J-��Ǩ9��'����T(��h�K[���Q���d�f�ܙ�N����q���e.,ηh���.pc�ԕN��������+�S����Ks�x�{�|��{���H�|����}Z�8 ��1~�@��޲)����	����ݵ����=84n�ݡ��%X�������ϝ��|9��c���c��+I���W'[ޅT����AB�afw���S vߩ3΅�#��;���w{z�yG�eL.k��h�z� �H�n<º����횞����Tx:�17��e���r����Y��/2A߁�������F�7��=�%�++��n�u�*���0\�+:8���E*!�K������pn�l��I,����,�j������E�����4��Lx<��f�u�Z�`A��x�ŉOa�d��,�����B0��]���͌:{љS['�zQC�����n��E��䣧��t�� mV��,�́�Y�G�_�w�y�Ku5H�[�q���UǺ��L4X����֞�2�jR�˚w��ק�}=B��/(����ٗQk�}?�27�P������p�����@�h�c��
�
E�Շ����mQ���Q�c0Dn���ϕĢ�WgE
��,ލcsW}d�J�6���(
I��cԈ7�E��:���� �7��d�Rw����ᄨc�����BR��|�{�@�����Gn�v[���;��E� �yS��ƍ��\zw��N��1(��xs���	����^��߄��Bi�٣�]}#��顲�B��z��R�?�In%-��:�s�^Vg-�������<Q�"�#�ҡu'���a�h#Zq>����mV$?���C�fܤ ��떍5Թ�ݎ��~�c����O��M^L��&=x�� T"�R��z֋������]9��@S�>x�s:5Ɯ�y���|>x�ғ�5)~�
D��P����[����K�W3y�6�ʄ��fa���WM��%N�}o|��yh�,��A�;V�Ia����J��+��<��R%��Yw]{���_Z ;�\��"_Ӝ��y~�Ɲ���c`a)��=\A��p63�����Y2�_�qU�zA�����W�~�r���rq*9��Pv�)i����&O�x��b���~���-˾`��ó����V(#��j�D�ꗝ�Bg)���.M�O(�Tg�}��� %4�O֍��cC2�+Ъ"J��MEC':}X���f<<][��&I-���J�凂��c��^���P�G��4߽ڢ��4I��-)��:`?�^�Y�ج�?��[3��KH���/(�G��JD�ky��	m憴����*%=I���#�mN��Ay���C��ҴA5�R�h���H8S�
Sʸ5^o�4[d¯��O�^�o����q�hb�ʳDе��,��f�	|�/-8��V��ԁ�6p�_m��K9N�Y��<��g�`	��v���NS�Q�$��p�T�烏]/��̈��ЈZ7��W����W؏�)��_9B�eo���LI��@2�i��cy����l�Ő��M�T�chjCW�۲ "؈����Bw��̀��S�YLS��ň������0eu���lUe5qO�R3�D6(۾��Di���D�=ʪf�޽��L�	7J�n,� ��g_�C�p ��3��tq��@�W�̆�k�̀�b�t�^�����㼰S�Pj�&�=6BVkvi
�fǊI>�瀈9y_z�]�j��`=�{ `s�{��
��x˱�����b0CE��R�q�F��A�~�����q��3Z�
�R\���J��Aҩ�;M����%�v�����sap`�H��2qZ���J��.��-���h����o�/���j���d(���cg�I-E�uo�F��\���G�]�ۖG��ISP��7&?Qt�4),a,��;S]h=��v1̓�<xQ{�P�mF�P�'������$�RX�뾮]+��鄾e�3�|f}��Ұ�7�ɿ<o���J���6��#K��K�dun���D���dh�3��X}B^�ٷ�sA{$��}$��= �YW�PFi�@]���X����a���2:Z�նi��k�c�_�nSjb�eǴʛ	�f��,�Zʤ_��v	��<�w
�
�5�*گz��㺎�.�'i:T����ٟ`�!��0����h9[��Y�r��Vo�+b�A8I���
b�1�N�����#����4j�ڈ��f����-� 1���*Ɲ�R�u����¨��a�oU���
���Dx<��?f!���y<7��[�H]ˮ`B^�� o����{�
P�z;,���ӵ�pe�"���?�G�,o?~h�:��5JEj��θѦL��f��>Id����d�:�ğ(����I�Kx?ܠu�M�6Fh} 1�o���E-j�!؋��v�`7�����0���ӵ&!F�ۦ{�pPG�ƤcN
E$Ȕ�����^S�M�g�z�TJ�ϓ�D�	�Gm!�`#�?f��3T��Oѭ�>!P\2����m��ݤ�ސ_��<��KߵJ%����I��	�����<�Y���<��>�"F�� -�S�^uf؍:��R������gt�x��U.*�UoJxݖY��M3��	���[�%G�=nߨih��oC[23�Z��W�$no��"�w+�e�	���2u��MQ�bwG�rdh�h��;�kb�)B��5�,}}x����O����8~����Qf�Wj��خ�*"�?���i/'��S��� k>X�M��|�℟��t�-c��(0���`�`Pw{������z=�f��8�e����F�x�c(�G���Ŧ;W����3'y����\8��T��Ӯt��F��������LN��E��}�/Zt헼�φ^#;eч/܏�.��=~d4�������Ԑ{�XL�����Lŕ�W��M��$����y&����HЂ3BJ����|�H�tG{?��L��F��49�ca�9}m8��z:�.7����jJc��5���A��&ІZd&/Hx"�R8���}�b�5���z��kޣ9 XT��&�\>5��TF��|Gi�EA���c{8$�|�O���;e�|}�ԉ�oOбJnHY/�>�phvRX*btr1�ך�/P�Ei��g z+&� ��Qk��`�L�d?����t���n�Kc���ՙ��4��i͠-0�.����D���0]R�+�$��g��A:׳6���&�)}�
���7G�(����G�D����B�����a��\Wˌ��c���)��=�[��7���U��� ��+����!�v6�4��;���fu9�3����rk��H��)���pN��y�5���!GHʅ��,�	o��S�tS���J�����ͼ�Sޖ�&��o4(�4��?#!�*0�޶���7�4:H_�����Ϭ��T��kt,��Y;���kc�`�䃧t���G��w���*�����i��+So��ڂ!�Q��2�����HC�H�0,Q:v#c3�h�����q�Z��f/�P�e��:�XA:pzJz4+Hɩt�9\�)A2�j(��p�z3�ﺠO��40l�K�@�ߪ����ٗ�`y�lY$ŷ�[������9��`��Kz���$` ���mT��|�n�����!Qp���M��N�9�1k���~�7	��`�������3\�K���^�e[w����Q�B�8B�*k���&���i&���j��O�C('����=������T��Y/��9=��M������I�.%��3�ou��N
�YT-��	A�*x�`�	>Nxt��H�bC�̧�́�nd���9����2z7����)i]�'�m����y�/�l�V��h>/wKA.}�cȟ�M_b�vL��i$�\�L_ģ���:��ˠ�i�jhkIOx�3Mq�4�c�;V��
��B�R���>�JN`��Wإ�����r�����mS�y�� ���xF*��� ��S=l���,�+~�u"@;������rka�1
�Չ��IG<�elIղ�q��{yY�;3b���Ja�D�D�����漢Ї�}���V���_�>gtFxq����L*��7��.k��}��<���B���t�߭О�x�H�x���sC�i�t7���XYnO2-i�Vzԇ)�9��X8&X�z�>˷�6��O �C���ҝ�m[��+<~E�9����B'�#��#�Ҧ�RHESD�sh��Q9���m$�J��N)4����.�[d{���$L��x�.��צ��3�'���E��kN�%O��?n)yF�Y �I65Wr��R�(W�_ah��X��v��|����.?5��*&V�)�DL����Osb4�f3��r�����yr���䈅�S�����|���á��2� ����֓���9>��U�v���+u#�J	��&���3�za�l?4A�������Լ&ŕ�IXˠ���&����t�C�����F0~��E�_��.(��g�(�/U���F���s�!o�g�M1�VO���&��z�[ �t�	���r��!\.�1�J����;ݣ�X��͟�&�w:ۮ^]@�k�K�e�8P�V?8��`� 4��[�j�R|��#5���v���(�^)�|�D�h�rG�Fj�qq,{0鿕l�������Չ,�I6�=M�㱥�j��1ψ3X� �����*&�,�ۊdרԎ!����;�aG�{���|���@Ma�,�NUƻˉ�".�@,�?=H\��?�:����Y���|̐x��3	��E���O��f��=>�,+���CŌ�Js6G����'X�)��dZ	7iz�ܗ���)j��]Ϙ=����@��Q7Jr)w�h��4��U9�n$����K/�uoP�D+������E�e�S/ߏ���jEA�@^���K�Ƃ��Han��,��(d7̷L'oʅߡD��=M%k.'�r��%���4#w
ف�TX��<�9qnz����_��g�;S�ך�{D�0�_�9E_�o�w�r_�<V�Pt��qƲ�v׽��n����7��mO���7�Up��lή�W5�"A�TI@�������M�j�GTڣ�ng䘊�TI�a��[� \��}������β����z41O����D�v]�ѷ�f��Hp�7mi�f�����)����3os�����Ft���I._}�Qg��SR��~a���}c���q����'��6��c��/~n�˱I��p����Q���-���Ⱥ�1�]gb%��M�τ)f:�q�>��#85_O���aݕ��Ģq�C˫��D|h�νE�*���w�'�*H�zppX_jG��hQ9:]EAx(ҵ����훯�������z�.��kR�K��1�tž���G�_��^l�]�7�c�����^��c�)sv]�1�?��9�/c�8<xX�+?�p����Knf��Β%6���p?�q����J-������44g�n0*�B���uP�Di�"�Ē��=v�>r"C�O5X_�z=%��M�ݿ�i�m��lg����}d�?X��:�X:��*XZ�Dw���ܝ�>� s|��#�c��w�S]��Sg��=/��Z���,\��u���H>��}�ҿ����@KǜL�(����������\WU��@�
X/<��O�w�9�@���4��f%�>�g������*�&�]�OЮy�',�fv�S�p�i���ռ��t�n��k�g|l��{>��~O�n�0����s�@�vi��$��K�� ����P\�/�2�q���}�FA��?p�e��nm1���%_R�D�,(�@+_v�rDť°ӛY��B��$"|I7 �$���%CZ�H��s`�_yȘ1G���7cO���inW��Ck�v`d �'.)j�H�P��o�����g��{ꨍ���%��W���+L�/��Rx�^Hy�{�ɰ��7�5�qf��^�m������7,~���êų��5�%3���e*��iN_6����o��{��'��J�o�Z�O����J[�BZRg����Lj(f[fj����4n �S��5�w1n�\tS�kJP�7*L�t��E�&��rI4��.���p<u��Eڿ�ޯ<����X��=�-��#r��Ej�t���x��t�iV1������wR��{��|����a�N%H��v�6���������
�Be¨�>�����6
��} .�?n��_��
I��؟N&���{X�Q���E4�����()Ň�������խI|����ï+M��X	�B��k�������ݧ�q�+�p՛D
Cy��[u� c�jh��1�m1!Hb�+^�A�9�#"�"�1�� ��"�o=־����4`��ܘ���%�
�,�1�n1�Ђ����W���k�$E f��Le��6���.��6�>8M^�J �M5��Սn:���x��<��1�+6|1�i��g5�邸�LH�iwxr�9<���Ι�4�]ӹq҇x��8\n�8����^-=ܜ�����������	w��;(�b��%f̥��>~�l�I?dW�5C~�z��������K�Y`k
�&Jo��.�^⚱ӥ������(kw���w�v�ݠ�B(���٧����˭����/���G��Ry���?%���i���ǯ]s�q�[	{�����Hvj8\ω)]�V���:7e�!�(��1-��r�3����v"���5���Ϝ�q��{��v g2p'L���р�q/�0�8=�`��jRR�wS�q9#/\��0�zљY���ad$��9���>*l�ӈ}a����EU['P�����a@~`�ߒ�>$n�$A�E�aZ�TL5�-�����x	^�:|\�h:և�)j.Ki�x,pg!��;��46P����
LZ�ծ�?�(���Mn����>BT���S��/�^)�����R���]FP�}ı[��:�3�>1����3g����x���O�Ԭ��=�)�.�Vc�!0S'9S���¥�h�`�eX���������O+"���s�G䨩�F�]��b#$�#��f��6�0�+��@�\[���2'��=Q�k]'M���pV���7�Q��}��!D����>�p_�?yMl*r���6C���<��qɥ�ò�\z�5�l|��X�v���w�Z�J��I�( 0dئ�h�_[�^���=Y�θ��Jk��֥t3���p�Iu]�r:�8!JG-�l�����Gi�Y�u�1��H5�{��k"�DAj���
RO�3�gTb���'���_���HPj---�)82��l�O��yi�u��č�_2��%����Lb�����V�#��})�ٚ�3����?�`�ldfÒ�}Qz����FI��Y:^w��x�	�
����^:�\� 
p���D%��{�SH�WO�aG�n4���s<�xv�4aH@+��;]��Ԅ�bm'�(�4w���_!� �dϲn xu*Y��,x�b�(����o��F:��t��d�e���i6��1 �k�S��D�ٟl���w�|ߗ|���`QH�n+J)���s?"W�<���6��jб��g���1��D2�R��*�%��Q�Nl���D���u�f%f5otV�Bf@�N���?�8�>Z�t�3~�O�Q�%!��aͶ���8'�b�Fl+`��O�A��E��x�.@̗���A�.)-0S��x�ҝ1��'�j��p3e_��K�����l�&zP�p�{�(2k�8�����md6h���+������a�7���k�-]Z�	qCQ%$V�3Z��a���KiEyQ}�\ ݩ\���G�
�ﻮ Q�q>�j)����I��%��]&��?�ݽ�R9ܗ��n驨����/|� �����ck�@�K�$���Ct��\N+�]v��j��`��V�3V{��'D\���9%1�<֪�����\܍�V=AZ<������0")-�b�Z���'k�v��(�9B�R C�W���wjud`l��t���������)�Q��r�5�P33s��V�<�iP�#N�RK�8d��R����}��23����F���;��MZ%e�S�2��D��,����:�W��יZ�m�`t�2�s�[��	��_L׈��J5��&�u+��xuD�F%��\1\c:�ͳHBNM��*"� �����fW�BS�D8��e$�*#�e��^8:nYok8t}�;��t����H��O�%������������֝r�s�n��������4�J�����d1W�pG��B_�����������cc�<���	7����C%e��[	�&@�gHuQ-Sʒq��I~��cr�0@�雈2[�O)�����>x[��mUc��Ѹ.�tyK�$d�N�#��S�=�HC�􁤯U�l+��Ϭ��w�,��~vd����WnK��+D�H?��p�������]��.]9��$V�GF�@̋qK}(�h���ڽ��a�&�$c���!}���Jh�vP��pq�_�Q�c��#�.�BJU�z{�9I��/����~� R`w������3�(�v�Yi+w7M�z�^�'���?�i�֑�hOrڡ�Z�2?�GF"f��[�3ym���x�6��4����|ta�ii���.�p⧘h(�R.�P���]o T�
�bc��y��JK�T�EE~#�*an+��3�ZEwE���t�������ǔ �����  ��@��Od-���쫿��*�ƬxJ(��`�F�k=��eQW$��U���4�>R���6�V� 
	��'��Y�'���Ė6��ݼ���f���ɥ���uk���FW�$`��8�Q�+a�<yKR�6�^�b>R��sVק�Ɔ4��v+�٢Q���� vH��h�.�M�hqt3�Ȩ
C�v~>��ɩ�w�x�.j�`��u�&�(<�5cN��g����t������,���bI7"��M�]g���ύ�qe�tp�@�A�A�������M111�A"O.��Ř13��Y��� lt���b\b��Nڸdt����ʕB"��e>�R����~}�owi[j���=��ņv$�~*�ޗ���(���"�GW�RπVhIUt���� ��h�c���Y<Bw�L�_:��_PQ}߀�8ۇ�"�_���gk��kI'Z4"Yd˨)?������&���]���(�yC���	��?�����c_J6|����IkpHk�,Oᑈ�6����=�A1Wƅ�u��[�SS�p݂��C��fܿ	^0�fFF"L���T)m#:MD����g��p�G������жԧX_k1��?S\T� fxf���f�����$���0��C��}r�mv�^�8�%Lnܼ.G��N���T�V�x�C92Ǿ�W_�X~��PW�k���'ŵ辋V|9��t�o��~�qU���P�Q�I}�s�����.8�AO3�B)1B��K$AE��E(9��t�SrYn�{�e���D�AW��Gl�͌\e ��B2��Fi��I�,8Cb�ܪ��s�)�vN��� A�/��#���+#֟vZ7è�%Î��t�k��_���S�w�.L��w�W���N�|�6��Ҏ�o�-� \l��!��O��Mf�;��e��(��-�_>@)�3_�=2S�X{��*A�BeIC���l�E�G���e>�2�h�誯}�H$�vhl��n����[J��e������%%��6��@�Zc� CT1��v�zaG��Y��4���y���l �ǏiC�3�UeR����0UQ�! 1f�`������Wm�馔�(Gqu2�6�I���R�� 7RmY �Ę>�6G̨�e�)�@����`\��j%c��s?��nXm//�3�?�x�O�z?��~H��䍴'�$���@��m� �|���SQ���G�3���2Ẳ.7¾�X��D��|(���2Dsx1�к��۳��i����������S�ƌ����|F�/ng�O���'��;tn����ri�vg�bK�Rv,����R�ƥ%�V�_��G�7b��ڒ�����J^{�h����Z[�pggg�G�͒�s�G\{M4Ȭ�+�J�+a����i���h��J��mk����;E��T�Q%򙒼�������y��y�SR@⦄����(�w'��Dv>�~�Ʃ�q+c���z�g&�<z߾sV���&�)g���"s�7��l��2�@��
���#�,��������2!���]�6�^�'*�q��o����R�h��H-��f��o}�ى��ux���A:�; ���(ϙ,��f���T�&Ѯ��V�����]��y��1��g�Gr�Ŭ��IM�<b���k=5�tL������r� ��e�x��Ǒ���������{LW��"�J���(�1
!�7���Z],*s�k*��u�����o������S*GQ��R|H���D�G��\� A�1�����8�ʭsaA�qb�������Kގ��������O�0����g��v��:ìz #��V{'E����[g�O��V	�U�7�c�_EP��:~C ~�MЕ��AӸtk�W�}�.-�%=dfڔ��T����s�I�MGpXD٭���6<��/�Q�<:m�;�?�w�?���g^P�Sy���x��)��q��Vj���V^*7X��X%��2x�8�#��RǦ�G+^=_j��;>­�]s�L��:8x� �Kz=�s��$#+�6ڧP���&�����	��;�M]ο�����[�ڮW}�ǳ��GY�C���;ir���Gz�DX�3�
��cE�;��jp� q��G#G��q�D�!���iK��baYTU@~.�v�-"4�N��#���"�:w�U��e
�|}tK�ɢa��4��B��/i,�+	�N����>��(<��cß��G�9�*j�%�7�☠a�Y]0�ۧ�W(+�|"��h�"e\���%�<5ʈObGS�nFm�I"�sm���,��U� i��0=�6��;�����V�Hd��K�>�~�D�\�d��@R�M�3�0N���.��.�<�zE8�R��4�Z^��u�ςn�A��չ��2�O�-AV#�f0bf*�P�ͫɺ�Cr|:Č>�L`Q0��>�
����E�Q����].Bo*�!Ƥ���k��ҳ�C�	��u�Y7D@g�@��^�G_�t�VWH��x�M1���0��.)�R_LG�~�!�#�Ό�c�0R���^���� P������ m��Adj���WgĠ��m0,�ɬa�����-_S�p�%��
Z�T�1����ﶧ0��CQlCO��+IN�βxi�t���+#��M~W&'��t0H7h���;s�80;2�7���P�4<exh�%a�@ŉ1.�^�ӡ-��g����u�*'������4�>@��=\z
Y�i�]PJ�����%T�R�۱�an&jy��K�g�n����I��]�C���@�|�μ| ߴ8q�-��A8l[��}���x)���$	D�YI��$�����ӂȮ��~q�@�G6���ٞxX����G��gÛ�jҰ�j�0Ϯ?ZB���N�s���XekO؏���cݗ�(:}��ee5�KT���?K�{�V��^�Bx4�z{Z7��~3�B��64�s�d��3x�{�+�lCֳ��מD���a�	��N�+g��������t�.���� yA���騅��Ò��yV,˽߶�Ї�d���j_9QF ���m����152 ���T\1m�3>�\@��u�L^QL=#tN��3�E�{'��N*�x���SM ����u�����������Կ�ࣀ��}��������:d��"f��Z-�A.R�f���=���A0���&��z�}~��X(c�����6�()�v[-�k��W�{��B�Ԟ��~�p�'�T�|>���c����bj�RYC[�+K�5A�����*Ѿ#����d���B�玺��}3P��tܐi���T�Tf<��:�n3�7�[ܟ��n��ۮ7W���Q����
 ��}X�%���B�Se-.緩����C@����]/!�{��݋d���?T{��4I�>wC��P�6���Y��ɉ�f�IU��"��ֺ�5�s֊}�>��d�g���ɠ��~��L�`��]S������� ��}+���stF81�0M'Z,y�^7Y!��ͫoك���U�Vd��mg�����}����g���muh�|z�F��!K�'FG6�aFޏ���&�E��]��hY����9��&3��=�j�]?E6�0���oP�B���+ڏ�)�Uߍ�Cn3Vo�D���{�d�*�a*M��mc1`�����A�A�k��*������2�}��=P�}�s�i���pzC��,�q��֮��9���w�Uύ���Y,l��� ���V\K��R��n�)���8ЀX��`� ]%b��/^��)L[t������"��Uu���x9���WM�Fe�A8̽��uᝰ�7�!J�Վ�/��u�+ܿ;�#E)��-�w
:��CbЕ"$V��h�K�R�<�>.�7���[ݷ�)3G�ϬJ\��S���/W��� ��Ru���AjO&�}`?Vt���̦bհe[�qoR�?���1�0V� ��9�B��ތ��*)�5�n��'
M�\R�N���ee�Χ��lH��Q?s��7���1�n�����r<�u�!�A%�>�[AR�>����wT�����Y�����csN���7<�&0�;N���#7�.��A�m�ft�{�3�����?�	b���h�v�bϮ�4��#�`���;�����q52D)�>�H�D]C���`Ʋez����}�^�G�<w���_¨��{ъ���Q��W8|g�~�!Qx�U����v��q��A�dҎ�=�÷�9��֫j�{� �!絴�pI�C� 猀=�j_�*�/"�O`	oU
����X�����ݎz��z��7�/4�4'�񴌦�q~Z�mG��N���k����`����&�;�2��&|��Qmn�x��eD	�1
�)�5"o�1^He���WO$�����<U�dOC�I/�2:s������~S³M��i���6{�y�LgyD�C�b���F�ލu9k��
�y�1����F���i�)�4=���?;�qY`��y3��8S��VT�P�����[yVi��s�VN����ГR�R�o���S�;(���#� ?a���!�s�y�,�a�E�a_4�8�*�|¿KX��y�Q3�ͩ�7��h�43�ۓ2��d=��3+Bш����DWe�����|;�P6�j�-�����kvf^�|��s��G!_+e�/��F�ۻ�9��[
�gԢn�_�������a�~���~	�g�K�jS'���b)%3l������_vk��J�L�����Nr-�.�̘������@�Z� }�؂�V��Oh���sHʰ��v5�z<��;�gmU�E��G��b��u���SS��� ��|`็���j������R�p)Q��|�s;+�6O�m�X�ͳN�B��^[T�4��J)K�(���:�J���j�8JF��M��*�~g�'��X���ۄt��=�࢕�����7�B�*��AW�F��N�K:h��y$11���q��Al�T��'���?Q*�#�lX�jm�b��|h�:�PD\ègs.�J�Ԑ��]8RCn��l��@=."����~'����Sx<9�P\��	0��\{yG�JJ�޼k)"dB�#q������e��ot�rH�uZ^>!�O�}�wy)z��L(��O���&U��(N {�y��S_��KN�>���~]|w���p<G��6
	�4k!gٝ�
��:�����$M��0��T[C���D��f�^v$'$s3���|ߎ�RNu�Y��ۚ�Y�pSi��PH���O���!`���}����_x0�w�.��u��ذ�n+
�<�����#J�A@�#f�U�+�3f�t @����싨^�1�j��LM���	_�8[lL
�|t�4���E�͈�El����^����/���,��Ǫ^���Q������n��:o��^dJ�B�Y./Jh��/��e�VE-�����V48�9�(��\�% �Oe'&�Af2������3yR�΃�bP�	<��㡁*���m�<+w����BYKelq2ᷤ���	��T��oN�覰��+��%;���hV�(̋h�gx�tmv"}8%I��� 2%��$�&�T�g�~���:V<�T�����"��15�ei<�-2.��{|����`�(m5xFĸ��}�'JS��|M��cr2��P�s{�MΟլ�^s��	����B8�<�%PF�����W���_r��:>e�����@/�"b�8�~�ѡ%9��OpY��Wj~6�>�+B�r�EVEi{X�駅��XZ�}zd_�>XT�%
�$�ק]�p ��H*��(KD��f���ܣ�F����K�GL�aD������o%�<#���|��r�`\��S�,B2˒=Z�F�[���PUu�"�,���Ę2�V2��`K����Ӯ�.%�8RL��"3Pox�]qˊ�9D����C&]���T�w>PB�r�k�B, ��F��p0��������wR]w�1�Lf���5Z�xxp�]_��OW�%��^��ʤd�G���Ȅ���l2ugȒ�o��2<�\��|�Pi��#�Q��4�sX/�3Ɗ��RH��@f��;=�>��K�:��^�����f\5���!)��C֣��qJ��9�6��OPB�N�l3�����jYc��6�f��o c��QC�%
��!�6�	�����+�ۑ��9BQ`�~�{��1mF�+	/P��v��ͽ,�ewA(�����	��qY=%��(��r%#����s[M�o=hlX���'�If�J��v�.W	�(;�Eh���h�ʧ��ρ}:��^����o�Z	�K'�&'�]��M��wgh�E[������1�����j#�dr�S��V�J�bb毦%i���J��o���|C#kz�)cQyt7�����>�&�֍�/�	r&���f���3�|Yo�b����fh����m����}_�]X���<<�Gw���==^T]Z���wb�50e�,T\�!���ʃ�O�ɉ���+��+MƂ�0��������|Z'��
��=8'��������»�(��w��X�A٪vIߜ�4��I!1uO���� �\~��o�I�7@j�(�{������5�U�<��K�ߒS4���!�i I�C�
��E��8ixT=nI$4<N�q�,!p>IE�p�faڸn��t��y��S��U�-�{{U�O̬��-�h�5=�*CE��k�V-{J�e��.��rK��c��-X�(�o���O�И�j)"��D�-3h�ʐZ\��B��h��k���<�w�WY�7�λt^���j�w\�ST?�u���.�RD����k�5��Jk��vnd��1*skG2���E��99e���u�\�);�=��c�v!�o��0�>�O߽��B����=��Z��W]<ͷȟ���E�<��T>�Hnd���ֿ���z`�.s�)�x�*�SR�Acx]�j��jN��.ί�.돞��e�h�>%���7��F%ꥨ�0��q�?|����ީ���b̕�x��n9�z#0���^�%O:���K��������������:�߅����wsV����)�/�Ⱦ�X������i���j��N�H} ��)`��,{�%��d�?�8Q�c�-Lr��h���Zm-�S�׷�X�?9`uk[��������}�v��z i�����p�Et�T��=FcU�Ց�[�1���NS���▯�$6�I��Z������K�箢�
�o��C�<��#$�ӰCz��]P�]��_ಛO�b:��n�'5}���G��	J��pU��'r�+]F�F�B ���K��C�,��1>�΍���ݝ4G;�K������h\z4�:4�F�g�z������G��3�u�����y�K�L����ExBF�;kii	�Օ+Bl��7������:��PX&�ݓ��W������;��k��X~K�.Đ�=����ųd/b_����>2����b���s����H����vՍqe�T�d����O�)Aqk%��̭���8>�Z��#w�N�Zm��q,����A�ȍ�e�:��	as����ߞ�{C���fAS�������7��	F��~Z�?�,Nג=�~�=qN�:���o{!⮺ȑ�|�eN_�|*�p�f%$����F:�įN4���=S�DϚ�/����0ځ�W��09Tr�Z��ġ��X���?
j���֪�ݜ{��el�6M���'�~6>[�s�-8�`z�@���F	GO��]VJya�/\�����H�H���L��p'�I,��^��������8���a㛺+k�nc۶m�wlul�6wl����f�v�6���1����j�D�ZK�?2s%>�ˡ�	���T��,lԻHCJ(��k\��(Z��Ab���v��g��0�纑uҵyi�e����fi�� 4�	^� >��'2uA���n��
sv����i�s���_�a�`�ES�AOz4!*VJ�C=59D X %ݍ5��Ā���/%_Z��.0ij bN��=X�5�;o�}��ޘ�܉���E�D^�7�[a���6��m�4x�`���E���kW�i8[��+9ao2�#i�3U��"�E���B3�DΤ�DK�)��A�NHN� �/$nis��%SLǆ�Q4����fJҿ��\s%05:��x�\��D����C���^쏴+0�Ej�� �QPGg�̉p>�.J����iV��[���0�W���J1#0'����tԖhy �~m��#1�UQ['X�·}t���J���PJ��&W��Q>��^����n|�؄�teln��}Z֬�ϓK:}��� ?��aW�mv��F�p�~�I�w��_����C/\��� V�H~<0��.4yy�Bٲ��jC&�ߍ�����@.�Ad�QM�<�%�j)���&��Ϳ)�d�q�������������!�J~�F[�����Dy�o�N2��:8N����J>O{'�NhY��&j��Ѹ�N��N��rqA�ozL,�V�!�Ǻ��ǆ}��5EFT Y$'�_loVxsW�>��]���rP�h��q~��e6|~�(�҉3��������73�{�ӭe��7H��E�~�َ�J.+"	��f� @��QE.�B����az��@���Q�rl�4ֶ7�١E$1�` _n1����b8�)�x�'�c�BȉR*̏��GQ8v�뇮�`K����]`{�p���eK�K0��%O��_�z�?\�{g�[!��{���t��,���C�Q�o!�E�h����E����~���%������2�bAb���<fs��D�h3�be�]P�=f؆�m��Su=�#�_���{�#�7(����;±};�q<s��-���h��=���⤊�ܰ��V�P1"�KB!_�В��t��3����v�p�D�d0Nd�&���`���=�f�����Xp���$iC�ݘ���XPU��N���}W}u�?�&�F���?i�^7��	/�OD��Vu�e%�'U�5���"('ӋmwAb����� &&'Yo#p=o�,�0��B�޾�����ZM���*�]��Q�KQ��t�s�FkN"�_v��3�`�����0�t�`�0��Ɠ����,��"��!@�.����fQ�v����\I)�1���"d�z��N�; g7}�soKjE�y8FMX���T֌$�_IJ�Q�'^r��jt�A�@��?[	7��ܠ�8�e�dq�A�=/�xO���������m �v5�c��{-!��8���*�JJR���+��(}��c�A5%��W��kQA�Ҕ`R%�o���e�Ɓ�}�0�������v��S����� JS;B^�/C�>�eƲ����i���s�C��n���X>3C;�����?�مH}+*�-����[LN��:�2�Ar-�G�M���@YE%x���x� �p�z���5�/�W�D<�Ҙ�L��_�~�I�4�Tq�'I��a�"�Gʓ�R�����
)���7��;��nd:YC!���7�Q Dm�q[��۹2�+�~�����1�g�^��z��Fp�+��9�3<�D]y�f�e���"��sy
��J<���<��������PZ�	�li���æ��6 �eB6��9��7<�?}�FpYp�M�	�۽##{r��&peɤ1q[�&�a����
[L���ܽ}k�Uy���<vX�q��=1Tb������1���h�
��:�/<z�Gs"�ㅐtl����X��&&y6��	(t�P�l��;���Z���h����;���jrw�Y=���H�s�#Bh舧$,�+����)����cE��8�PMeĭ������d�*���k�T��4L�ʡ�;w$�d��!'�$��a(����E�k� /f��s����~tU���Q_u_�$��#bxs�K�h��đ<o�K�ϋڲ����������>�WV��$f�gxD��۫���uL�1��Q±��T��(�0��倆I�3�� Bd[d�:#!J�������E�g���4՛L6_ʨ��������
�Q�]y�v��)*��4t�\Y�A���$�_�H��a6x
���m�Ԭ�@���s�F��2�SҦ@Z�Ud���B�'Y-trG��n9�o���8A��v�ZڛnJ^����o��DGu(�)�_�
����3��%P����@ ���-�Ɨ����N���b}N�g8����+�s��anΣY,�H�rx	9dd�Y�x�nߪq�kc��N�pUyʑE{z�?%��:��uyr�mW��h]��7�#�[���v�� ������$t��U��>�#�B}N.�?����"ⷽ�G�r��ʃ�۞�fSy����K'��ذ�V��
�	��>���K�0��^�V�z�敻	v$��3@s����T#�{���c_��V���̻3���ܠ����3� ��K��T�E�.���ʂ$Q}nn�F2������et����{"�\ѡ#�D�P1�5���>R-�
�j�h�!3�~���8�>��	UE�/����@Z�R����9S�����.O��R,��k�]g���;�3<�}��֢�J8p�A��py�U��TO�q��r��?����d���a�o��Y?�����e)��Z|%�4oHݩ���X)��N���7�á.r��"r�U�1�`Vs������8T8!J��Ug,i�1��0�a捍�����9o�p��h,�Ll�s�yV��3l�P�Ƙ�$cr��_�|�>���jpZ��kX�	5l�����zX����q���/+�~�S��0"�T$p7���7��qQ��r�ˉ�""����[��ݺ۪�Z}j(���M�3jf�`i�c�-�Z}��T%_0@+!�+5�b<4�7<I�����������3b�(&U�DN�!H7yc�&�¹G9��Tb�v�"����[qq��p�S��v��+�G��f��I�O k3��'8RULpO���% ��Ќ���V#V�'If����<Of��w��-�K:;Ks8�p�rÐS�Z��=�IE��lCL��D����^�|s0��97uޅ����$GfEה.�kV���0�4��D�!�4(�*��]Jv��1-8��LV�.�w�ˆC�-���P�q&�*Kгc�����_���&�Lzwz������������[��#������E��B��������D�`E�l=E��+#���k�&oF�\�:�+��A�_�CѼ��j��p�"�=�s�HG��Iu����ᴥ9��V�3	��D�y�w��:���Ԥ��*-�4>.���o�H��@�)C+���)EG�P[�J��Ŷ2�����ktֱ��T��*|�B-	�:���$I��BJ
�RG�Ir=qM�}��x�Gte���+� b�.b�vSU�uu�k>�^{d:c��g�w�e*��4B A�b�52���z�!�Fq��j���?�V�+�a7���gjy��6,���U;Zp�{���;���8G���
	O�T"-��K0D��Ad0�O�B�@E�6Ei���i�H0V�u�:�i�a	�af[�&�4�/�Z~�G��?	4y8�`�u�E)8f�dQq�]糉�0
�*��f'|�r�����#~�O���+(0�NB��0��N%���0��z7  ��>bZN���P�"K�

P?��H䂳@�L� n��Ômvu�ߩߊR!�i@)����	��\V�����ua!��J0������ԁ6o�"j/nMUut�Ȧo̖d��Q�|�����\��0x e��&w�WM�`�+������рϋd8�>i\,f�K��!g�V��C^�Т�l�Nk6H�_���e�*M���cKR��U��lk�_e�V�_9�j1�cǎ�pλ�lk-���`!�H��&�X�g�ԓ���g!��`���F���؍f.R�~�6rf�tP-= �+�a�qKQů�G���_K�F���I4��n��\�-r;��'��[���o�`�w�z�x�gXT���K�m4�]|�x�7�y���Y�\H�29�T�1�d�9��L�ǖ^�|,ץtl`�p!��X�u��.7����9�X���~ـ��f�����t�Y���%0�4#�NM,���Cp|x�V��$?��5Ӓ�Y��� 3�C�7>��ܠ�$)6�����/,3|�bnP��;�Pt�E�5�h��wy=��S�Ւd���v�!v\��e�6:V\Ie�}-J���̥��D�$*�q��E�#�!�A���!��DS}R�)E��	ۖ:�y2����EY��xi�G+Md�q۵TR�O~e^���u�v"1�a���ǽb`��DyE���a��=���k![#�f�IG��<���L ��<�>F��b
����n@q�a�}��Įa�?k|��:{�/�RQF��>H�35�[�G�l:��eJD��K6��	��c���e�uJ��I�A�5���pgU�3!�("#�x��Ce�p8/˖��9}��o��ܲ�}[ed������Z�k<�J;K�ş�������V�� h���\do�΍��x q���?= �I�`Q+������늎�׃po����� ƍ�1�Cÿ3�0@����@�h��A׼S�H�a�!�1��fy�ێ"7�v��ȵp��U��YT�i���8eE%�Ro�[�3f'�خc[:I�?g\5���z�I��ϫ;Hx)���)��[�Iy�IM�b��8 ����g��[�@;�I�l��(U��������H�`�P�B�`�ێ���;�af(g���Ks�	
N��Y*'��(C�26=�~*��=|M>y$:�+Znc+bQ���"Ec2�t�z1�h��Z̛��𞌚���cB6���C�����w��<�������G[��:���rm�v���X�ռTx8���UP�g��ױ��y=�״Â��j�\�8�[��]�.c�o�p�8�n�޻�F��T�K/Z�4j[M˵���i����.�}��ZJ_(��� BK)A|٘��nmS��֥F��H��vL	[(��_�$�z�ߟU.�7gTMn�:%���w�j��91����ʒU_�GGUiJ�e&��>�Ұ邧@?�Ö1��f��;���;1|gp������w,�@궼4,�T
r��F?K���38��k��U���؎��n�C�'Q���3<<ݸ(��۷����s`�L}��M�F�v�H[pƟK��5F=��/��.S�~���)U�nc�q�r�_fP@aRme��P���T�̑dˮ�Z�$6Cyq>hum���[�an(;N�|�Ԇfg ۶w'#��}B��?����I�1����ø����] ��3���}��ȳ��wr倀A� �R�-���2��<�>�'U�I3ncBm��W��4G�	*�U��L��##������5Y����j�Yr2t��e�i%=2~4Ē%�i�������JG��] �݈,��[������~o��Hc���<6q A��,H8�	��6UG�R�kJi��~lFk�Tgy6���k+昸?-%9`���+=�>�ԓ��
!Bw�.���AЛ��qe|���X��/U�^F��e�l��7��%�lL 7(�3@s��ƶ�(-rC��u�|Hw�\���`�/�a�]���!Mܬ�T6 .��L���鮷�X�t�|g)�sB�z�+xV��>�=e�Z{|b�Ĉ�$_���*|z��Gs�c�<#�����}>ʒ#��G? �S�ɷ���rY(�k��`��wr�B�M@ �}:��$󯖔a4~>��Q��u���*�F0�(���i�qM2m��F+D.�4+:r�G[���	篺:2�O��t�N��tc�5���[}U�E !�Va���ٍv#$e�g�Udbg�2Px9q'��m�H�����<�b��JW�~m�����s�p���D`�[�]�`c���T���
��V�)���g�7�#B �wJ5��|$yNPhP�̇U;����~��|!�����(������-�٪�F�|�go�YfX�oJڃ�E��"��;��x#2K�/X�r�~�P������;)�~�j�k�[K6DZ��Yf�6�)��tV8h��(O
�h��D":�Q2�Uuu�:*�`ܭ�A��1��1��_���Tf���z`�h\&F���he/|F�B�K�Y��#��k�=1k��X��O�I���K��O3��YO���J��n���hTk�Py�H����YƁr?�\�Jr�;�Ū-ߎfU����H(xM�I؎���DѢ D��r�m��B;�O������1���`�~X:\����Rԡ�<�% Kċ��֛@!r�����.w^Ne��MN�!�$�LL����[���;�Fۧ�wO����-���Ӕ	�$Z��7u6$:[�SbS68��\
|��ٻE�Y[a}(K�����/��3P}�9+��F�15T�#��k2*^-��E�����hD��z"g���*ͥ�����Gpɺ����D{�}���\.e A�逯�PNx�ڧP2�9�2�j"��+�����Ϝ����G*�l�S@)wE�6c�}E̤�]�!���D`g���������r����i����b�E�^{c:�=G�L1Su{$�"n��{���@�`��[�v;����	w6���<��f3V�#�s�!dc�	\Qtcu��*l- KȰ��ȋ[�6�{ɥv���՞��'��ʑq�2x�Ua����_��5��V6�N�qq�~��>#T=�	���%I�/jF�'�N�ۄ��-�����nly���tGO�m@ ���z��<�O7=�5�+��Q#�tyl���m�ݡ��dx��3��*8X�	�_�D�W
�p���lGҧ��R�̼�)v�۲J�-�b�F!���R8�A�J�R����F��1�E���_�X��\�@�⅌鞖�H��&��v)p�{���%�(K�n���#���my���u�͆�u�`@&*i ��F�˻d��lç�-����Zj�������
��կ�jRf^J��!�
G��*�c)��m���=Ġ�Nf'��<�7��a�Gm&m���?���·��V
�;�V�O�A��5��Q�qX��_��t?wN*
��p���϶u1K.��z\w,3�s	�48��)qI�eҺ!E&N�-O����td ��I�L�|�#@��9�� ����)����k�D4s�^����;���Y#���ѥhf�,�A ���J5�4��l�ƶ[cg+"�?�>Z���p*f5R�z�R��$�zd��_1��
,���c�,.k�M����4�}�2^�n�rds��u� ��Q�Bb��[y�Q>ǎ������u�a��y*��a\�a�9�F�Ф�2�}Z�ؕ����Bc�W�9����E�DRQ`�8b�_��*�'�
N(ɴ<��U�VͿu˻��*ʀ���twb�f#�cCaj�c�p_��m��ʶm-�Cyz۸��H���X[�Q&��]XE<<S�zx2h�L��խ��Ό15Te�kE����r*w���p��&S�0�^^�g��V�ہf� �s~of| �B�vF�z�������lu1����|��:�7X4����s/R��~�R7B#/�h͞;���4��!$`=ڌ�Kg�R���� �,#�	G	h��ZP�J���L��g��UI��7��m����ܸ��$U-_�J*H����"�r��~����w���`�\�{�t� l��|6�'g���>�w'\��7�J���ń\ܛEC]�!D�@��^ϯ�Z��('�n�?�	?��d>��Z,���>�p�!��M����`�0@��L�'i(	��'�OC�c/d� ^4$!r_m�h�`/�ލ~.��'�q�_�$���𫐎��k-��q5g.��^'����������R���y���>z�����d� 0�x֔���z��Vg���h���&���F��lvt���W
�d-�JH9L��Y�W�(�*Q/C�ȗ{�.�!^
o��w�)=���I�5�<W�<�*�4fv�n���� mC�����`ۖ�RF�G�1�Y�z�|/n*:5�_t���]��\�M/�gu�(�FN��������=696_� ����ӡQ��{su�a���w��Go��_s�/j2C��o��i��xI�FK��w��NF~, c�!h�f��JR�o1��;��|���|�4tP��"��k��$�PR:�!5iS��h(���O�ò���ȉ����ʁ��}e$xh�p���T-4�s{�w&%�/OU	gpN�,vpiLz{&T�?8 ��~8���o�k�43�"�F�=��`���[���8p�[V��p`rZXR�r�23b�E�t&6�lݚ�^lb��z�Z��
�<� |1ߢ�(p蠌)]8:�pR�"k �8 �I9[��}�6�{�S��d�x��f-�x��gU�əFh����n�mb�$��:�	��@Jq<���DWM��6G�`&z_s�3�^����K�y^ nP �^}zt?�"��G�m�����+�%XoN��h0�	&���N��Z6�jQ��Y9�s%�z��aß��Cם��ٰ��`�$E1�F�vב�&�N?��y�9�B��8Cf�"���d=eH5k�&@%?�{�&��ܻ�	W�ȅC����>\#/,n�Y}��R�2]�w�_��kM�v�-�S�=Q"�";4�K�6/=�T5C%M��G�͇��j"��\���<�l\&
�)��Y/m�^��-|q,j�m�"H��G V��*U���
�k�@p-��5W�;�3ؒ���6���	LKpS�/�^�}|�9V	���|�T����O�\�pHbV<t�,��C7�ۥ"��鬖��Ht�����T�6�yh����D��^1��h,�^�sB�<���L�C��=�Ŷ/9;5�:l������,06�̓��4��H����O=,E* i������<��d�d}7!z2��3�y�������,\��l	OK�/ǟY">?0���ly��MI�/<R��d���|$F��	��C���U�99�gFj�5��ITp\�����˚�
C��k8k�9.(��9u�m�YS��D~V&���SJm�2E^jڥ���� X��rXC' �av�+#j� x?����c!Z�s����jvz�v��֖2����4Z�Eò��u��d���?���
��� 5:��'�Dkc���z�I��2֌+���D�i��+�n�SM�����ܹכ�:�"������K$6/�9�/�}	�s��+��u��зJ�`ü7杬�c p.�	�A��6�OEU����5'�!�R7�7�ܥ�g4�.	�A�M؊ۮ��E4y"AK�n������]8\����QR �I�-!a*��G����R���_՜��lƝ+�m��j��<�|�Xl(vvvd����l�q�M����i2D��J�IB�W5��iE�\������e��YK� �xuq�x�6�E��l���2팩=�BF�7����",���]�������6�Y�2Q���(jk/��~D��z��IU���o��<�z~�R�-I���2U�ƍ6�BEE7|�3k�!��L>&�x~��g%�a��/v�C#�������"s���Ƌ���%��/��|��k�VzD�Y��p�P�����1�*�_�7����~Pk8vW�y#:���"�$�[e��Rh��#z�n�#)�{0
�X�k���y�p���f�ܴ�����K�"Xb/��*A5;bv&��L�w.`(����K��ɳLӽ�d�۠u+����rK��R�L���={,�fZ�38Sx��I}%�L~�1*�MP�3[o�$5?�?�ıA8ى�K8rsu��Hq�fx3\�EdF�po�f!�ϵ 뵁}��\��=�'�9 ������v��ˬ1��l,���E��5mNhѲ2+��v���)��?�=x��` ��Rۃ763�6��/��4��\�w�+m��ߚ��y�+*��͡�����]��j���6�
� b�I%�}����?"�2?:XƁm�/�ޚ��x�HoU������'U�`�Rt�����s��.�������Ag��4�.�'fO�)2u>U�r�dԗ��������	��V<�W@�cF��Ηx�(�ϻ����i��)�E�IB�8x�8pp�vcw}!�d��n��L��T�J��m�Us��|�HM�*�	L+����*��w� �R����L-uC;��J�v#-=���sqvg�1��ܸ�������ў��%���c�y@�d���댏8�{�hs|S����9�ΠI���Pک~���jD�V��t�~4'�)8�L��?>�J�v�q��5��!��Vo���x]��"�C�6{�y�tKy�\�ψ��[��Ϋϊ,_9���D��G�&�]��7S��W��\٪�.7h�1\/����{��D�������?t�@�0�O��N_K��ە',���S��EUv���o���Q]�1�M�jo(�(�����]}k������eoW����6�@	���K������gJ�fM�Q�*���� �+V-F�ڦ�E����7L���V�6�A�B�.^��N��D���dA�ϴ�b��!e-��{l�W!|\%���H��ù�����Wu��ǣ]�q�K�.�m#�U���M�N�՝��^/L���<T,3k���%� ���ϩ���N� �����Z.Ϗ�+�_YT@y���zBX�{�E��BR Uq;@�BW������:�Ds���?X����R����_+m�aX�F�X^�+[W�R�ȅ^�yY���F�E�Jxo߉�u��l�a���,z	��ݷZ��Ӎ=�ccT�X#1#�Qcj'^�@��PX�M�����#�	�� !}�%M�� ����iǂf�O
Rj��p���c���jf҇)^貅�g���'%�܋�|h.F�P2�89�)����!���;-oF���K4W�n�6WD����r��o��F*U�{�^v%A����Լ�Oʽf���xm3���y��#�@9����\��n���ڎ���݄�.� *0����/I"&7���}���n�L��&*�����/��:+ s��n���s�5���o�c��}ņO�"eK-���
�qQ=�`c\~�jZ��KL�R��M��;����*���+����sn�Q#C��sQu m��<N����W��jAGKأ�e�'(�H�U������̅�D�tr���IRDI ��*-ib�s;��`~F�	�YB����=�a�<Ű�>���b�J��0f��#�S�#(�ߍ(��A@�@��2!�ޮ�礢�Wr��m[�+u�b���������2hH��f�`,��(�37�\����]lU�&%��D���3�e����I�s���Ǿ�U������� �N֞����{+Z��-X�!����S�?�p�K��g�qj�5�3�	kP���o�� �ô}����h7L��Nh`氼y��`�����w+�g�%�iD�|���ru�X�I�97�e<5f+����K2F��?[[�$v��e}x��ŗ'U�i������6�
閒P>J��{Ҕ�$n��Y�_�2��۹�cyo�	�����\n�!���{��jzy�^bj
K���N�M�J��=��&�z��� ��S�%�&�bA)fvn�a�V�㴑�-:�ۙ�g!�v��ۛ����դk�~�1���ݴ�)7sV&��0�Vo1�~��}��GK� @���D]�I	�P�<����m��rÿŰq��f���A�!dƶ�� �y87(+5��خ��#�P����Q�欯�D���?��}��}�p����T��sZJ��r�%�1���pan1)�i�$(c��#�5M�Q'z$�#e����w�Ý�/�Ϗ�<�5mm�YTA���k_���y.sP8������������l�A�9��+|3�*�ƈ�߽򻎭�n 6(9�̂��A�k��{��m��S��t-���y�&�l���J2E0q��EH �ѯ�j%�x/h����r����P�����D�� 0���������kn���B�H͕�H4��&�ͮ种^$���$�_��Μl��cgX[�������͈Q�W�@Yq���L񵺝�#K2��v����~��ޥk{�d3����bͭ4��*��ɽ��k���������^��|�0��0�?3?������V_;�[�P0G�ow
�h�����uc�B��<���k^A2d2�(H�/80C.��E���ݬ�������y�Y�XZڈ����H8�� c,�0�,����*�7�e_�~ٽ�����������+Ĭ�SLcq��4��Z��B��ʼ�2�f.�A<6��`�`��d�9v��611�q�Qޕ���b}��Axã{�;W�2���r����ٳ�K?�E]�^U�?�f֓B��	���I����`��\K>J;�M��(Z4��Rb�{��1ύ*��H��vp)���rum��mW�^������Ox���&�4x@��"���RC�篶x�Z�]��"T����wB\_U:��e�	:�כ�Ź�@�Z�ۘ�h�{���Aw�uv��֦cM�xR���vG?\�l�"/��� Zޡ'�C04�7u��f���Xo)����BCV�� U&��(��{���jل�lGeY+(�DH�MH 	�sK�ueP"�G��k�����G6���;�ֲ�������Y���)�O�R��]����&>���d��������|�����H2���Z�B1�'(b|���*o�Va�b��sB�/��>dF1��>d=���m���<� ��/��D]�|`�3y�{C�q��zv�-uP���5�.��#��\?�9/�/v����p������2��],7�Q��}�$^�q��M�[}���;	ɨ�J+�j�&�	���r�G��D��l��k�rf���+:j��XB����ӰSGԓM�45�.Lﻼ٦�C*��,�v����� 
a�MT�����oi��W���M��XQM��%,�j^r��5���Z�;��b6:p)z���fGyM������B��[h�x?4�`=ٕ�Q�}��ove{��{�C q��"�ӟȧ������sfƘ���޳H�ϗ�B�!�\��u�����S�[�^���<� ܹN�o#�7��{9+��Ov�O�J��F'7*'��+�����*�	��d����6D�N4ϒ��!"����1fF`��p��U�>ApXj��{&F������V=G;%��(`}� �4?�;�5W��Q���G>2��XTƟ=i�)p����]0BP:�\Y��o�Ã�^A����ڡ�"���r��j����V��ԋ��
6���o�8�����;+���O��[�j�{��+��u��cL����.���]>����$�T�^�UV��m���l� ).������&f`�P��>h���
�Fl�����ƈ��Ͼ{8��7(�Nt$�@k�-���A�5��-͞p��d��������ߠe����h�t2�����m ��j�)
bi��kѵ��������JOt�,� �b�����G��LD�?���ZC��5�"Ӥ0��D���I$�Z�L�R ��p�8�9-�Q��O�q�\����Ӫɞ�� �u8�Y�zZ��+���xi��>Q��z���-�u����A��6���p[랯��7�f}��5�b,�[�Ȱ�é�����U����Ӆv ��Au+���?�ЧoSĀ(��_��t~8�ȇhT8(#J���ˤ��f�(�3�� f��)I�D!�՘�?��6�52�Ff1D��5�O�����+��
�	�8�g��,����Ă��E���=��!
�,�m�$�ΗV�sY5j�6t�=GO�"��HA��VB��r,>����w6 �*~Ц/ą�����TP�t�r;����0��`��מNT���rQ��X�p�����(�
;�c���*Bny0&Q����ׯ,w�i�~��]��U;�b�9EC�{�H����'�rOQX�_�=X��'/���
�*O&�O���U�$"��Tl��q��r���=�H��DS|U��t�-����x��5�A,�C���^���q���Y�8���Kbq��6�E��1��j�;�=�uT����OM4t��� ��̡�"�,!nd�
��Q�ܽY��oC'AE��[NИ����^�{��
:.;v���0eݯ�)E�_������8x�s'�M�B�o/Nx*�Y�Y5.�E�p�����W��rkey)uؿ������� �G!��,G��%��ԡ�n�E��.�[@@����Df����t��0`����5�t?W����"ߎ��n@��fu��;��\a�`5[G��:Հ�
��=H��\R�赞#��aƠ��@����/������F�e!��}\mw�l�q��R�L��B��%/��8��T� �T�i,)�5j.���v�Ҥ�����-L㈂@2<��Ϣ���X��p={�W0���Ћ�����^J�;攓Vr����qe�`?��$�w��bJ�{�]!���30�:@S�b{�5��N�p��^�g���2�f����to�믙SNٽ�����L�OoՕ��N�MS��g^ף?F)!u�X+�?���oxL$���=�I�n#B[,\w@p�BP̖�*S17�N�VD\-��7^�ؠu������38����#&OWL�\�EV�����σ��ʲ�6���v�H�h�({�6ܑ�c�j߽k�PCt�]��Y>Wy'iZ�8��6}?T$�H?�dZ�$L�(�Verǳ�p*PB7��0�\^h�B�X���jD�NC�,1R"וu�5]e5��:���������W��q���!����ݓ:Ŵ�8���#2��E���-{=�*ض�(��b��,އ��n���E�նZU�o8�d������n��Lȯt���N�G�~�xh?�����|��x~��V��Ғ�G���D�^/~v�ĜZV%Juv��--��^H��4�M��X�dY	�
)���A�q���=�iPxw�^����1�є�K����-m�om�� ��X�d��(qe��.T�Oci+�G�f�M��Td�����uC�K5��	a�j�]�Ժ���}�u���%��>���mB#�[7��&q<
�5��'�0}��+<���o{�������9��$�1�5��}Ύ������ pI�rNyj��C ��cO	�Y�eh���aEY�F;!`����Dc������<��hb��ß��}U���#���ۙ��)3�A�ǙWN���*<����LW���!�%K����2�����Ɛ�Q�^�H��
�H�8���ϥ�~K�LR�}��b�*�}����H3�nd�U�6=	m�D�SG޻zEh	V	&�F?�Y�7��K�|
mU=o�V}m��P�~<�b��9�_���a�8@��c�5M��߸ʺ��\�P;��4B��B��2�o�q��J�ލ��%cE��$�ˊm3��q�o�u�;�մ,]Cg�[�z��5x!���Rѵ}:N��A��;~������|}����A�jv����/|0Js�	 (����I���|��D뫀�'�82�&�6[���z\�U�]�/�����M��{]_щ� դD"S�&ҏ'V'��rXo�8��
�`��0�=/W)�+t�f�ZܥDK��7o��Ɖ@>w��!kܟ�e
����qhGz�@[l�lq!�n.��Un��\�^���V�NJ�w��|1_+��`�}B�}��{w�v�L �q5ޑ~������cs����X�������x�_�s)Rj�'TI��_���:--~�х����s�f�˟�#Ȱ�*��3� qo�"��W�o"?s���p�~�Y�!�t��Ӄ�y*�dF���M�H�z?s���/���������p����Hf8���ud��#Y�l�Ȉ���dIV٣lQ�q�qQ֑u�p��^G���>���ϳ������Ck		�59I�ͩ?�͏��	֜'�	�<��wFcEQ��T��]W}��V��y�d�D��x�������J���/��3v�v�������R��r�G�2�y�jb�Dni9���jf���'zw�LD�o1�~<t���$V�C�oT{&y' �3V����΋��d�i;�=ى!x��S�(Yl@�O��ǯ4-.�r��T�+�5�?T����X��W����1��|IU��;���\F�\3����K�l,zZ��Z�vU�;�ޛK�H�r��w}4G�7b5]�w?�*���H��G#�
5�}��BF�]ܾ.[z�ʠ�rL��S�\���G}�A���qM<�7�]W�5�o:��SY��4�����z|�؀:G6Y'I�Knl(�����~��:y��*q�q��UG�Ķ���[2(S3
Ѵ��M�(K��7�i����m�[.(��+	�P��/�� �OG?�6rs�ŵ�6./K��V�д�aŹ�Յ��? **j������jyYM�'���m��95PR��gj�wG�t~������|1�+�<��{~���³��ĺ���8C ���|�gx���坙�f!�"`��/�y�8:��P�+���Jb��1��T���bȹ�O�.�y���w����zo�nmQ�W7�����3G8�)��ӈ��f��H��{K��N��Ƴd[���k��k���F������_3 ����ET�cX�������@)Ŝ��b����_>RD�ϒ�0�C���ZYO����l�{�ә�ٔ�6u���e$���<b�&�^s�Y;�飨284�@<MQKg��|��3�=��*w�p���ĭ�q��5�f}`�T2n�0<$'G�_�|p� �ݩL�?��gin�p||�s��H�W����R�ҭ��wE߃��q�L2�����,�g���y��܄٤����o�%jM�ʗ�ثpq��7���C2"\eO�1),���45sB����0�5�uzx�^2z裛n�ʫ��V�l)�n^6(6�pK5���t����C���mL9H�~����dJ��9�i~�1�Q�g:�E��.���'�iQ��Ɵ,~���"�tѦp5�%�%�9����Yi)RD��u
<^�}e��w<��(��<�=[>�=�hW��`"��3���Jp���w�a��d���5n�U������bC���$�F�D8�;'�;mԍ:��'�H�nܴA�t�z�+NEp�(��4��C�Merq�8%��F�fA�i��yQ�|�ԋ���ƚL�<.��W~��b7��R�`s����6�N��9���Q��*L8x�0a��
i$R[󥤊����2B�h����#���2m�JJs�LD�bL�-����������D���G��S�r+Pn6���Q�\))d]�%#^=�1�k>}������	s�^!R�M��LwuZ'vj!��M���(��a=�I��w�K�4��վ+�ԣ�6(����ah��/an����<Va<�Y�u栴�����Ň�h��$f������'מT����],�)֝�I��;

E�ɫ�c�;�`d�8dӗh4=����5� ��w��].O��w{�l���0�s�3#.��K��e�t�����g �"�p��	��֣g���S���SҪV��y<%S�㲛�����)8˾��ЍWX8���o�ئJ��w'w_�`�Ҋ�Τ�JO�:-�ܤZ2�H�8@�EO�}'8��B�cT�1��ii9�@Ê$趯��gN��.��J�������W���JiVvgrj��F�O��h��/��qO���u�!m�Z?��ԚNޥ�g��0�>8����K��6o������k���<�=ˮ;�W�!�c����Z�����}��ӀS�;��݊����e�X��,�U�Ƒ�FY=��eF{s'[��8�IAY������ʹ�����b��w��ů3�
ˁ} v�B���,�n�:ci��_;S�ر��Ԫs�T�8�:���=N�ÏK细�%����u��b^���2�Ĉ���_EԺCW�O@������V��kL����O('�l$���`��P�`�A�|���+O�R�g��� �".?���NF�lT��7`��S �5��2?]�Dq�Y����rJZ}9� �*Ȩ�
꼸��F�D���ɭU���>1�ں��@(5�װ���?p�-5{}Ȋ��m &t�
\	�Q
9!#`֝��u�K�%�	WGš{��_�R3��2��������B��Iɷ�:?�w�查W�3h����T���;���q~�{��p*�����*��o��j�/�HQj�"���E�ȍFF��5�T�ķ���\o
�-�AE-,��$�#Ra���v�� `Uު�(T5����Lc�̐�1������+9��xs*�zQ������$�#�kj	�k6�A�-���~G�p��v�c-���鏻UA�sH�u���rQ^\}&E:5]<mQ��+0��ȭ�:_/'�J���JG�B�ׯ�;;��r�'��~=�,J�G��-���D�V	�i��y<�>:�-)j��;kxx1�"R�y��;v�)řy˓���5� �||)�j{�z�{ԓ��{��iR�O/f�������j&�?V�Y���k��-�ZT� 0�������V:�~��w{�ACMf�sB*0�b�R�1��O���,��^3�p��/цu0g�	���k^5;����Lۈwޫ/�:Q ����ǎBձ�1��/�E���)�*(Oӓ�� �N�j+!w�l�f��Nӡc�;1)l,ط�I��C���ЎO$�N��s�p��[���N(��������;��I�3X����:mf/��!A�!�3M�P"+��������{�L�-G�|�	_$��ϸ�V9;v����&VRX�R/7��}K�⁛b��O�ʗ��kVy�bF���M�x�Y���w'v�yx/�7�ɲל=)��������~�B6��c%[�.j�V3]�]�?�]tpǭ��W7=k}���~/V.ךxV��Ũ}�� ��ϳ��w�k����������p�_���C�s�@u�R�X�/UK{���od�Pz+/��&."������y�G�4�2���&~���NM��p{|j$�� R"�}P�݄+��Q��(t�^�Q~B%�+�v����g�����S/l/ �B�s�A�_��/+�ޫL�6H�&��f�^��f�w�EސVMK-�	����������p_:��[/r4��.�֍�����ra�!@��O��L�Ƿmj�,!�ct���<���NZ�e.}�"�|��Ƥt��~6�hoxj핮N��*ɭ�4�<���d+a�2x&����UyL����ْ�W�)zh�p�6��%����߿��<Ș���g�^�c��\�N�����PW�Q`�$�t�{r��U)/���ڼ�L��,z���yJ��f��3yڬ�x+�Ib�̍�?7�+n�D�wNfׯ7��ޡ��Z���շH�XŸ@�.(��s�r�_T{b��[+��r"��?���	mr�sQB���k�z�Te�ݼI�x�c�����?|kf���������v��4f�͸�"�7}m��N��PK   �|�X'(�5W �@ /   images/4737cce6-ef6b-4e79-82eb-dab57378d86e.png��?���?��*�N�Y�"<)�J�q)��+�9/9�ͩ*������i��"����ls�a�9nc���~=���O�].��?���t�^o�wL�=  ��߿� 80 �<t�w'�#ĕ�c��]}�C�O�!�������[� ?v�{Z���n���<�{q�>}��B�
n���O�;+@^�?�5D� ���~Y"}�~J٤��@\�,�m��g�;�o��]Q|z� EC�J���2q�D,�۬>�Xk���i�_TO�h������T,��@7A�}½���_ؓx[+��3<�������9�X��,v'�W�K���R��2���W���&��0� ��ِ���MA��+@]A�3JY�`���=Ɲ][h�Fq�M�p	@�3�Y���>j{~����;D�oy��s��-��y�����'���������߷��o���۾�-' �o�����������Y�w���9� ��2H*T8jfVtðKݠm�촿�h�X$��p�Y}���03a�H910�aUv�;�bg�"�gC��wf;21�m�1��m��K���0vTss���t�bbf쒻����|��F��C_���\7�.�2�%+���Q���}�Ȫ��dVO���7Kj-ڲ�v�S�o �>� 6{H��@��|��k̰���D���Y�>%QO�Kߚ��;9�ܠ��ܯ:�E��g��"�4TfIW����^�m"�ck6?[��;���qz��Z򧹤w��� :(z��P�F�:�G[\�'#�vg�#jKKʸ��Z���W`zb��+A�쫯1�\~(�J>�T%c،��&��ݐ�N8����_�h�l~��}�BU6�2���|!�`�u�OЭ]mz�V��"�����"��ձߪ\nC#�M��E�`�,��OV��H<���dP��)�����t�ӕ����E����O�.9a�q���:�bug���(�B�xg	������T_1c`T���Wcɟ��jܺɉs4�7k@$W,y��.�h��<^R�Wo�!����|(��/]�{o5Hn7�ǔA����4�//�蜿���%��6̋�)�J�6��7�a�/(N�˻@��wмiL�~�[�SLi�$S��q.�b7�_*-���j��Z]8Dj�'�^����cRe8��_�=+ZS�N����X[��MuF$���I/`b���=�nboZ�A�z�����n����42�����3��9��5�^CQriJ�>t�֖�q崽�j����֞EsV��,�(��>�u�w�8�$1�L�sd_�s�3R0Ոn���������r�bZ� ]߅�3�i�w�?��,oީ�����R�Tb��4)�@�{��u�GvލZ��GL���^>~ڥ�|u��,���Oٜ��W��Ij�̈L/|^7)��d�̰^��҈�	���y���	��v`�_o4�}��;[zoå�\B��fk�4N.������s����Ы^k��nH~�p��"�!gb��T\�{�O�L��t�K�Iw�����Rdl�d��B�oR���e�m����D�����h�qC�����Ҽ1.�*�>Q�>��c�8�
9�#��DVB���o3�mI+��5
mT� �hR�2��a�L&|Bn��^;���nM��}hq�W�΍��s��*Ʊm^A��xy�ڐ���ã�_u}Syk7q�	KeΜ���mC1*"Sw�&���(VT��-��>E��EW�t��ԫ�M�ce�.6{I�H]�sl���9�עQH3Y���KϦ��*��.Vj��g:rb$f�~��	m�'9���S�Z�Բ�(��2�s�,����_l���I綧:�J�B(ra�����l�.��ɬ�h�������H�v��/	��´"�8
�u�O��A��3V��3� {����|i!A��WNp�Ah��0�"�����yC�Pʾ���U���.���ه1�9IU�-�v�_��|�ɑTwƥ�0���۸��Rh��љ�±g�ckt9��OE��Uֻ}c��M46#5�2�����s���3�wNp�d���}-g�'�w ~��+�_{���UZ���\�m�XiI�7�r�'b����d������Z��'�t����5B�:Q������ti�-ܧӔ��0 ����!�ݎ��#G��ǧQ��5$�KO.�/��ԣ�P#�Ẅ���1z��]�C�>Z� �c���	��J-�ʺiZ2�xT�����@�>��Ӫ@��$�Gكg��on.���;y���Օ|p\W���E7�R���>9&��j����)�ѩ}5�$^xF��J��
�P/H�����a�w���ͪ)�q���Ie�G�
�dq�]��2�CBv�f��?"������U_I8�ڳ���4�R��� �}A�;-4S��j��:��t��<H93�O~|�A���M*�&�s�@����"jq_E/��1+�_x8���T�S"L#�I*_Џf���;��T�d�MSҦѩc���I��hj&�#�~��L����C`tk�� >`db�7�x�2CE� n@�Eq!�@�`�8W�׻'�w%��Z��<�������vw�>�,ͷYd��P��}�hy���qSǐ7-IXg����� ������R$g���l�^�|�j�6"�Mi�$,d�å��r���\�ۻ+~F�B��M#����͉l�����,d�B�k�G�^�ɂh���]���Z����q�Hx�C������ګ��f��nC�?#�d�<s)N�2U�RX�g�lWz=!.��H�^a�ח��@O2�,�����:�6���\g~�	ix?��z���\b���6��.rRU�u��Y�t"s����ya�4�����H5O�)`m'��x�e���n��fF���%ڪ�������(�{�7���}�L󻠫�)
䘱��9J d徵ΦtNr:)�=�S��xBN�[�9��S���
B�L�6�٭���'3@fKe�0����?��_�1V��L�����j�!��#�b6�>!��9�i��������XO��c����/�~З���eb�nj�.�������ey�F.���_���+���H�8�-!~.��%�C������9]6lt1ьh��-��B�D�݇;u�\d��]��C`JN�Q������AY�X��q���S�Ry��֑=���$ ����#�o����T���F�T"��9������i̦r�5�uٱ�}7�}T*ВM�q�Șy����ـ����!\�S^��&�)p�´E�<�_8)�3�i��m���8\��{i18W�u�Ɓ�M�5M5/f�Y�a��~wr���;�s �Ҙ%��|��REټ�#9�W��㼪�?3+�2��z�d��#�-'�"^��������Ra�}Ϯ�j�>�w�hI���lB7����;�V��/$wv��=�>rRK�
s�3�	�宮�œE��,��k��x|����,�w&$�]�W2Z�׵dD���ywEwN��w�DX�aN)��F �*Tca��m�.�Y������]��I��$�}���=¬ _,�F����s��Yj�W�n�>R��LMϋW���=��MYP�B�|ٜp
�I&�I�z����039pp4b��2]o<��d�`�؞Тg~n~�����C�����j�Um�<��pk��;I-��͈ȹϱ���."��/�o,}�X��-���z��;��M��sQ�zl����T���I���m�by�hz��kqv�����<���e���%�0�'�^��BN��� ���5���@,�v��n.C����hf��Х���	a]a���Iޟ	e,EO9�b�`��)#b�]���7
f�.���}Fl�H))t�)2�.]���9櫻v1W��m)D�2��[dow �Yx|�vw>��^�>f_��]�ߙ^��s7>�va�'s�ŝ��{1�1�4�ЏuW*���$��L]�>J�@�~A|��)ז
׵��A�~�[�\� ��?)'5�̗�{4{h`!�1��^����m�	�{��AeX}1"�Š/�����[ooA)����}r��Ŝ�}p�i&A]�P�Ik�F�F�`k�����RXx�T���X�i�X���]�^д��k�1���s�����3�5�u%�T��u+B����a�V�x�m|*^�^�g%�_��K���vֽ_��aR������h�����y~$6 @����k��{�~�%^�xb�o�����V2c�����9�6M+tc̦,3���M�ww9����.���m+n̥��B`=Y��bĶN�[$��o��%s/���a-\HqJ���sS���(Xg��	q�F`.e�x�������@�"wܬB�m��|�.�Bv-�_,���~�z(�_���b�������č�Kގ-��:��'�C��P�J��D;�Y�ON��)}/@o�xQX��t5ؔ�P0��u�Y-8;�EN8�*�F������n�>��ó	��x��ƌ��srZ
uHX*WJ��:z6���K�g��ɵ#�V�ZI��喱
1
�ea�e��j���c���!߮ ��Q�����AD��!�����_ת
�G��R7�6��O��,����L>�i����^d)O�s.ډ��MJo�����gh�U���;"G��bi<��$*�2�E�N��ԤS��}��@��`Rv��%͑nR����9��chU-�5���{GWt�-�$'�=��"����ǜ�k=��Ij�ɢ� ��J�ވ�y�~��IY�[	��/2��R!|��4a��?�����+éO��x���Z�G��_^^ܣ��M� O;�r�Ơ�$�X��c�{ �N��M흌Ɋwhi����<��s��7��1o��~�����'��S����!���:���ئ��'�6�7YM�!�
 �F��F
��4���o��"x�Y3�"U�r����i�݉�oOن"u�c7��m�����H���*�A]SN��<�1vh�����)�=1�Tb�������������Y����v�֮�m�/��ɀk�������m����FП�c>+{		��UjV;/��sx�<�8v�V�
��d���/�Gl�*Z�C�|wがQT""�ioTMء�^��Q�;<<Ί������X���s�~�ǜ*y�~'7��N�d����Awm\��D��+周�e�ɉ��P�z��C�k�I���\U�V�Lu�~5$�K#Ex(�g�%.s�o����S���\�F�{|�cv�����n�^\�69Q᳦�54s�����1ƣ�9v�o�ho�ՔL��Ȕ��|TYZKl��Kd��J�WC�%wY����c<��ؐQ��;6�����o@GK�[ܩ��߉Lr��h�(J�!usD3�����s��?8~#yg��t���~��Z�̫49$��`��KŅ]X~�O��q���.�<L�V���,��ǹ�J�.�-���cvn|���������ƞD�����>W�E�YQ	�ח��y@�ƪ��D�����p^N.�z1Sbu���*���İ�U��:�K4��h�ac>���m�۟0�W���ZbGޯ �_�ym�#qÉ����X#�=wnb������e��M/���v	?h9�N�!���j�i���=�7_��cby�#7�5�џz�g�gy�95�dw��'����CJ�S�/ic�Ãe�� �]���8y0 б;ڄ��S���t��A�icK��O���V�*9]��曖0��q³��;uY��3f/�1!o ��V\�:�z�^S$���)x��Q����
�UL������|J��Y�����/��sVY5G����i�^��*sL�J�q+�f�\«�X�P�v�6D֯G*���!kI���\�Nl�SŖ�zΦ+�_%0�~����R7�&#�7�y�oN��t�n�=tp�x7[�N�C���h�j����F��Iק?�)ğ3b#��܁����W4����O���d�Tս~�2�s�g�p�7f��˱IY���f�^�N~�݃����./*�:44�)T���#�/�<�/y�'ܰԢ�� _y���i��#.�n�^�9;�F,{ȩ4�=�����.{I)������r�4��(CY���v��_�<(���/s���'F� ��ޟ?N�~��=8w���r�z����I׈�'X�6u�~�,%m|���sҜ�y;{w�X`��O_��bҁ��VY��>t�
��skŨ�f��tR�T�e����|���`���49��9���2�^�~�l���ˍՋ���ٷ�q����%/���w��R�~��Ϲ�z�T/mp�@��w�5j�~�y�%9���H�O�f���Q��و�P��T>r�7�����>0x��8�:?����r�&4Z}lI(��$6I��$��2р�|4�;��'mt6����'2�op��+Msg)��jՂ M|����	 ,|OS�1R8!@8�-/y�ߺt�7�'���-����I�;�.�OK�C�a�jw`R���vSM�DH�$ԑ'�o�vQ	�CN<�_��h�A{��A��XU�BsG�B��bHY�9�rh��.�����.G�b}��)�M����S�x.y��^1���*y���3�D�ڜ��9ިj��f۟g��鬻%�,�1 F�|��Xp�b�u����s�2���� t�������hB��8+�좀����y%�Z���.󿑀=�^�Cb��0�#"ě͋W	9���OT����� ݗR�{��")J1&�T]j�J�aþ�l�)?�?����V�i�ɦ�y<����'D�*�<a�d4���GAD����r�w��-Th(:�"����"���)�uu�ʁ��[��fM೔ӥ0����]?52��-�� x�u���������}��5_ͷ�hx(�����q��;�
�Q�\��	h%ۤ�(��m�����3՝���T���s������H��+��Nq��M����ˣ	m���G���(jE�gy;���7���'`�� D8z��)��cw*C*�5]Y0�|��r��-�9$��Ϙn�i�.2�
Q)��uv�(���\�Gh�紨l���o뀦�)4)�\�o]�r�@U�Nb��eZkr�(�{������!�?1|�{P���d������)���kdF���6.�H�lZ�����W	�����	9x��. ŴD���?�봀��T%א�,ƆX�����ZC��4R��}冑���ť5,��Su:97!
B�hA-nQSיMAs�ugjlO���:h>�<�*���à��C~c�X�錄�X���O��X/���_]�L�3U|���|R����Dt��Ӱ� ��g���������˲m-���f�u_�=�i�ꋖ.���
Q�	+B����s��J��~�n�-���;��r�p�m;1�'��D;3��jEt.n�� �����/_��_�������3'���(���EK��$��í,�����@��z���fQ0�_��>���?��0*��<"z�� <[�'Q��^h��w�c�~(�L�����\T��{����~�a��N�f�Z�2DO�֗�RXJ���N4�R6x��"�e��Զь_+�9�,/���}����E�Ǽ��m?�n�q�ո=��!�a�}��6 ��=���fч'�M��j+�P+O�j/)4�|��`�4��U�!C�����6�C���ôl��LCO�h��]������Ԝ4����6Zo��L�b"K,�/�k����Ł���
3���_d5t���fD�(��6q� �+�`���ol�^U����~�>O &�/y�ϵ�w�V�u�y�t�nο�ؖs�Mg�T^�Rӌ�NR�����BBdiZ��Ρ�$�q׳�[M�'���C�ۦg�����Aҏ �ҋܗZ����K,�*y�f�syM]�
\������R{(�{U�ȅ��Ë+B�R��*=�ۀ�O�A��'�(q�z'z,3��!u�Q&Xp����c�����$��s��n¾t��O?�_Ij��p���`�v�j8���1#�bWL�}�oK�7L*:.O �o�׬������$t����7$L{y�=86}�v�bb[�RK�KK���+����];��sssWh �����;
�Zv�Q[_��_Nj7����R[���7:p�*�#	�I�k��&��]S^��2���:%��9��[��J��H2�^�iVONd��1����u٣�FB6}NU�Fmp�!YKTmbQ�1T,����iX���%*�Ol�_W9�an'S��A�4�P)��7��Zx�1O;3�G+4ޠ�?�ɹ��H9��s�1��2~jkl{Z95j\�O)���p{qj���
]
Ny^��d��*����z,��9���?��~����{�Wݥc����8#���Ps��՚߽&:q �jwz<R ��Y�qW������˷]q]gQ	���9&O ��o6�5R��|���Q۩k�/>E�e_��'2'��}΢�<��8S���7�f_�,��sW�Lb�F�ȥ�z��MHc�#�:"=� �����q1�����X`@�&hǩe�V�Qҽ�钷j�K"�fI/���� O����hT5T����>�9��^O
e��r��K )ó�ьMqz�EP�v� G� S3�(�q#�̞+U���9
��}j[Om�7��Y�(3�v�{��ot^��;9*�q��C���G��������ĕ=B�z)?e6,��X�Z����JS�[I�M(�`�J�ɭ��^����DU6II���0����w���_�c.:��Q� ��L�"пbc���ȑ5�w��>�1�X�*����c�ڃ���WEed����ࣗ3NO(=�F+��\q�bV�d�~܃�e���RѠyc��H��L��V��P�^�wi^#�����m��̻~�@!G��PO�٢�N��{�~6yY*?)P<V�Ut�va|*a-v�S��a�
;m��i��3x���}�n3CX�Y.mX}�Zoc��/kd��Z�|8��􇴯�s	M;w��?�W~�����������Ww�v��%����Ň���|
?Q{miz���'�Ow�o�y!6�t^�|6_���lߧr=���B�����9o?��g�8ROդ9M��I����Q���g� 3M�֏p��� ���A���s�7�m�0m��L�0T��CA?�rp�|�d����)iTg�Ͻ�	���r@��슢��SMXN��<B#,>Q�ˆKp��\�L�-K���G��d�1�$���q���ieaj% ��]j�o�-�Q[���K ���
�9^$�h��2ΌF��������_O;t�6������� ����	�>�*����6~pD�܇`�`�=��ƕƅ��28�J�p�!G� CI�������s��ǐ�zY�?�<n
�A���:�z���|,_��Ӽ-��#�@���>��@�m��o�.:rH�G=F_]���p:g돐�+x##|�a�^˖�X6W�
nFo'o���[9�ƭa�u1�vWX~ڰ��  �k]	���r����mz�79_����N�k�j�	w�� #mTO��ZȜLH��(N|V�Q��dr�����9�~�����AaxM%-��[B~t�A��y<l�P!����Ƀxл?n�  ��yc��!,�!��ȩ�N�����I��_���RW>g�8�*��K	=���>�8�㈱�i5Gٟ�dv.�n�2�Ȟ*��zO�G���\`��W�K!��[6m����,��K�v`���]Qȣ'd�yq)G*��.��.Łjұ���A�)X������'bku'�"�c�2؝
�o@����[$���Ƭ�7�-�+���.s���"<�u�����XI~�v�mI�1Dn
,��^���^H�{��]Q�D� �����
$�{���݅�K\ V����BqRp���i���B��5�	�s�!F`+�{]��	�7�(�{4���H��7���Xb�����xf̽�yfο^��OAV
H�ʁ�a���P�0]�z*�=��2�""�}}�8�Z��㴑J퐐�E*���e*�֟}aegg'�{�.~����V�ڿH����+��7S�,��5s��@S'U��L��ը�0ݸ���o�?����$�
4Ʋ���С�'hz:c�����C���Y�RifT�b�v�Ȧú�~"��<�ӊ��b=�D��B6�1Q��Ŏ4{��I��	�����E��>>���M�M��V� �W�\��O}�r����/�>(�RW{�3�����x+*!141�e�����7fR���5�^��kuL\\xlͮ�LN R͗|��N9\X�`�#µ	���Ek��THQi��=)�8�6_9y7��f��r�>�g#����?g��3;��i<ox�ܮ�������XH�����cu��H�������� �-��_��}�j0�q k߲L����9�\\��^��?G�6�zL@`(�%uV$C�>z�Q:���Ij�=A��DƆ���"3EJ\p^]g���^_�'5A_�Uu"�-Жg�·�@�;��>��<$s+y�	t������sg2Uй8���=F�m���|#��ǎ��rV���My��|�i/��	@�����^��,l;�A0_�Ryg��v@ߡ~��u~��8�u�b��%���/�}�.6c���{X\]�X�K�����U��\Ͽ����?�)f�1�����^��NR� qE��G�����<Xg����].���N=R���!ja��o*�e�R*L��������[�rj�=�P�[TT�)x�|?Ԑ�^�?D���(��Sg`�ǉ?��j� ��ʨ�!���[m��m��_��׻!�O��ǧg�C=��3�(��o�m��l��
�I&&�H�#�i<t���'��Ŵ�0	�W��c"�$H!.��<v��|��0v��6!�����������.�E��}o����g`Y��i5غ+�G��0�e{��?X��Բe銃��a	����x#gA8�%��0)��#�dO����S �p>&�恄���	�-0c>n~��� �[Ӂx��7���&߅��Co�m��,���#�2��)2�ou����l�qy�m�Ѕ���O�<�-��Β���+�ˌ ��EQ�#4x}�|E>ux�D�s�'em��F���:���*��l~�Kl���P��(����ɪOOW�>*�<�(��'#�/xIQ?߈"��G+9�_�}=�j���-����
^�����ȼ6��f�bx1,�J:�(��[�S���h��X���Ƚ�F�_��7Cu�	��̧�����e�}^�����JjRUb#�'��� =�Xz�v�,)�Bح��s7{&�W�C�}*Z��aצ��2$j��ޱ7�E���� �����p_H�v]�ZcN� 7`d���!z�{����8�޷@s����k�?Y������������|�ʤ�o�|�?u�W^8���O4����3�o9_��h��,%��j~A��s�G4YF�,;���[�_d�7P���
�.����PRR��N��Ø��/_��j�?HB{���BK���!��:%iQk�W�^w��.f�ܲ�Bim^ck�{�?v��*dD��|Hn�A{rkg��TÀ3�"&
�S�3oV�4�4�`�XX����ٶ�Q,��C$��8mg���$���؍!� P�7q
.�eK}�񣖢��$	$(��'}0|�7�����{��l�o1�q����j��#�;}��"PT1�)ͱR d���A�f�N�ɰK�=�G����Ğ�P�5"�:��=YS\]=�^5Ը��˕c�!��b0Z��*¤��7�)u�Ch�<j^Jr�-��C���T7�����Kd�(��Z룇�������ۿϩ���զ�g�\�ޭ�%��g8͊��#�M|U����&p?�wu���CZSէ�,Ｖ8�.~�r�i� �дy��эO��?���R[*�=�	�/�l�]F���m����z�`���ʶ
p���5�fW9������'������*���ڍ��~�0Z"�A������JG����Ɲ�rj�ֶ�|�/y�Jiٚ��*�0�2i���
tS�92*�Zz���ohŴ`mxI�,�=J���mQ%+d��L�^��#
��N.��.w&80ŲyU��ɘ�G4��W�@�e�h�T�?�O3�WN�;W=X�|�.���)_hX��,7w�H۰�!%����H�tC���ߢџ��ME�q��S��gK,�4n�K��v�D�[IcJ'��={e߳Ί���Y���r2�0�|����E�?Q�,|h�l������G<��SF�+�D`x��	�*�&�0���4��+Ф#���h��D/{�x�	o��>4S�w�{�<��v6������7=����&<*.*�}*�Φ��20RL6_�x�Wɇ�_��.bP�uV�Fj͸�k�`�SJ�g����[}}�f[����t�U�������r�2�v���O/��
`桩��'	7��S�h�J�GD)�L���K�e��g�1%|w�mN��u0��l�i�y
�V���t<~e�˛�
n/�vJBRC�I$R�o$`19�^]���o�T4��d~x}��ώӻ�< @c& ����%�BXt(:��7�T%/k�2k�a	��@��J�
�]���!���AK�Ű����\�B[z�!��o
WUSU(������zT�TИ��� ;���UL�"�jb2,��ШQ0k�\���)�m�e?��6�a��I��B����ꋇ�R���J�}��НL�����+��ywd^>l�	��~?��uJ	Ainv�ܝ�.2� �x��t�t�uɍ!oւY�!�<�
�X���PB���*�K�V��"���^m�i���'y udȢ�0L%�Q�^����Ⱨ�6[��عǨռ8��3|�3c��zN4:�
�ߘ=`��h�D��܆tSW��{Wc�s�!Ý���ȗ� *����h�I=鬋���dK�%��~��{ı��%��www������(��z��n�&J}���Fh��l]p��uʕ�w�Ԟ��T&I�����?��v=�}�iYf�>xB���se��To�/Y��Z��ļ�dMZ1�-��p;Y�?�A�1�k�I^n�ɕ�vW=�[��*P��wX#:An����.�t�Ʋ�<7cE���wynv6�_�E�FZw������?�e�p�p݂Ka��)S:�gF�r��ᓘp{R��=�6��u?w����.���i?G�{��{N��)�����FM�������_���\�Ǝ4�Dߔ*�:~e&�0M�K,i��y�m�du���só���>Z=$}�lKy�ְ��N��6p���6�w���J[037�#��s�civ���(qK�U�A�ST�.����*X$�P)�7o�{��n�eh6OĮW趒�+ӌ��oT?����U+�nL�~���$I�Q��鷀����;�s�?���\��lY�49xk�W��---[�`���U�-c�8��F���3>�tujsR���ր��Xy)�	��Ϡ=G��ո cy�Q�שd����R<o��ϽR#=�����t����[�Gm5��VVZ�ɗ�Y��P��;���`j�����;���(��g���&�h�3NM-s{�f-,\P3r�LQYi??)˦	N<z�P��tg D����
!f+��fR�O����)��pc��EK�k�Xf��&��1Fx��Hoↆ�V�4�@ �G{�2|_�n��ȥ#K�&��+ޮ"�ޮ���R�����Z:O�ڂ4�Z�:�[��roI������{�n��v�`r��m�����PR��vwX	�@y\���9�k�4

"���l�ձ���ּ�6`�K��-����
S�U8�2A�9�7e�sH�q5���p��@J�Y?� J�F��e�իW����`F���S?H��t���$�ݾ�ߴ�:0��ѵ��C�nD���ɐ�kw�����o�q���J�@�_*�����U̱+���Z�A���4\�K�(U�"��=hg�%a<��>M��@Q%���U��'�$�XϮN:'�hΏ��>�2�kg����}�e`3B?��]���Z�b�����GWA-�U����BK^)
m�z�~��)�2f-"���x��<N��	��|}}Kȡ<&:Dg�y=�
\�����q�����~l�}�Q�V�^o�a�j��� ]���jJIf����f��������pf�17�pV���F4����w��CPڹf��:�HJ3A��`s2%���X;5���h���C�vGs���FDR���@�֗^E�g�
W��w���4X;[.��wp�&���lc]����a�YF���,����XҌF��Dť�p@��}�ۢ�dd6��M��I2k�~ސ�B%��3B��4\�.�]e���
\~_�XF:�P��#����YV�)z�%��k�a޼�U�ߣ�04z9n�wG+���+�����%���rؗ|O�?�r����Pl}�})�BC�zZJ˺�q�R�dg�Zw������c+�R��|���f/���U��C�yn�`Q���Kz��@��H�MH�OQ����3�P�{j�X�������b�:��߃���nR=:8ܴ�2-F�����Ԩ�W�"�E�"��]�/!U�y/�\���U}����'�u�X�Z�\�|@Y�vh-~�_�x���
0�-|
��qJ�o���E�w$Q��i����R�ȯu��M�_Y�ʭ6ɽ;Oge�۶�B��RQM�5SʴvN�ph���!��vm���_c;�/C��j������8�G`�<
�򱃧ԑd�6iL��,uYb��B'��\�VZ����T�@x83�b�jkj>� ,�a��~Vc�f�7/�a[�WK�|�����V���=������TC��iÏ#G�ի�"#�q�+���9��C*����>��}@�J����!S�%7b�̾2A��S�];�Py�~��|V �gY�~�Q�S-��� ܢ���ȑ�{�4}޲�I����Qr�Қ�?L�9����̀
�%�;�e,�_|�N�2X��߻ #���6��pP��}(B��4@�������h�VeS���h����z'�i^��`��v�O����*�H��Kaas_RC��SZ[�9��.���Y��:wR��T_�L��E[��C� ��A�X���@4�a�
���`n���U�6�=O�=-1W?����î��^��6=
f�حK����-..?�i�eA�;�"�7(�ÊA�*��Wx��� 5��8;�t���{�qur�9-}�q�_ݧ��N	ol:*~k�􇰡-|�"�ţ���� ؃W�Y���rj���j e8�o�˧_s�Q�ي����n��+l�	�n�ƹb�F������'k��Ƥ�W�s:$�I��'��l`�`U�Vvl1��6�^��"$R��az���CXicꈦ�j|/{��#x?1�4��l%Y�eETh�eʳ�,��n
�y������uK�H`h���cjf����l�#�9X��J0�3;����KS�3��Ōeo���e�k-g(g�,@Qd�c6C��.��0Wp���P8X
^ t�5� Q�'?_��q��q��]p/��N~���}�y���z3k�AB��e�gw9Ws�|��g`aI��MtD�m�fj�� 3n�F��:�Q�m�`��5s���t�cu�'��?���q-|��W����͝����VI4fH�$�������St{Rl.GC�o�(p�QP0���4�Ԥ�w/u�YPūqovӑ�-��ձ�N�X;0TJ��X���0Ib>�`�a:�d�����-�N�����L���H�fM�����9�/J3�a��`^�I�=�N��y��P�����;�i�Z��2jӱ�H�O������`-�S�؆<�Q<�z'��q�~�~�wƏךT�֡�O��K-r��e���3�z]�� 㼈�O�ѩ/0�O���ơ���U�]J��!���ٗ�N�U�!A�?F�+Qs��=��j�8q�/���	~1�v��l��QZ;�[�Sc��L~�# �>�LK,\�0����A��TIH4H��&V�����S�3!���j@�W�����kN������G�/V_�?iK"���[��غ���}m;��c�c�)� 7}��ф�kRhƏ��%���@E��M�cZB��b�A�j#������-����j�
:ʚ�YL��O�$���ǖ�j�ۅw�mvH9�٥��v���%�}����*y���)*��r�q��[|��"�8���ݏa���h��s�	}���N�Ci�{�]�Z3�K5��mz���L���d*��]���ׂw;�������#Fd�7����g��,�=.<���+ok�j
ߴV;�`S�dV�V�6�.��z�x��[����`������*�n櫶L��>����<�����/濎j���RX�
Y�Ⱦ�w���m�
kZ㦻�C�ST��9���H���K�k���e��Q����N�<�}
Y$����S]��J?�NO��t�PԷL)[�Y��L����1��qM���8)��%R��))"�"���0:�Q�K@0�FKI�1F7�a0ꋯ���x���������{��~�$��"]im��H]#Rj�~���^��mk�2L�I3���q�G�T�L��=��CD����hM*��>_[>(`����Ŋ��HCOc<��F�7��Wu�Wq9h)IGj��:�Y�)�!Ă�rS���MvV�~��Q��tM�%�=W�Rg�����������5�V�x}�{XMܞ���B�z\2æj`���=�;%����IxV�[@5+��Kj�K? �\/8����I��!z�1���M������}�=Ǝ=����bjS͋샺mD�T������38��P���/뻳qR^�k��L���tS��p'��P���/� �޹�7b�~oi�"��/'&\���0 Ǖ�G���%���շ����ʗX�^j4�4`���ĻV��f��ӇWJ&��z@���1�G�1Q��t!�Vg��>sV�����k�D;Ƕ���]�MYh{N��)_q��6|r�E(w	�k�'%�*���v����N:��\�dLg�g�O��>ϗYLQ-�V��%�œ��8��e�͢���.���{n���;eʻt���m�= j*�cfw��SH氛�几�����.-ޔ\Ej�"M�Z}�R,��5��nsX�$V�$˷4����yz*PO��L�X-��{-�&�x_e�QB�@�ȇ�f	��m���;�h'�:�)�X��=�=R��|��gH���C���7��/�F)u�2M?cbZti�\»��m���e����ˀ�I��ȫ�|� -�6��׾�R =����1��ߜ3v��mB�ކ���\���3�i�Fm��n��=��7"� ����8��y>�Ɓ��Y4��t*�{x��8�����c�g����4��U�"��j��iT��s6�R�8
�q]�	��U-�.A�����5���C�r���=�}dI��zP�������U�͍�`�ۦY}-�j�G��7rO6�{plνl�}y�� �:)X��sr-�r-A*� T�rf<� ����!k��U�-� �>��I�G$8��s7�)�ڎ�+vi�g�w��Q�����Q?�R�?�;�Î��4�*;/�>�}zt�n{�%�tySFEBok˗�l�e
d�^aI���y����(��Aӯ]�b߷��2�>�`���7�?9�OӶ��l+�Z5X���خ��m7}�S�TMX�v]7�,[���b�ٯ�w�R��)�����n����ڟ�#*�,
IIМz�����U�$q:u��,�F�Ļ b��5I�'��:��!���v���4�3\ϷZ\m�I�Ȭ���I��q\�]���U|�r�Lw��J�?9T�!~��a�;�׉��	Nr&{Df�d���.��v;!��{�	=�f63�c�P��(�kDy3,��G�1���m�d��)�j�X�̛h7�?`B�[��&��.zze��~˷%!Yf򋷐i�8 C�{���U�E��K�7����W'��]�^lPFz����q��d���H�+�A9ی�w�5Y�-��]n�P��m<��W��-#L����2F7��#s�o"�+ey�x0Q��7i ������m	g����״�8�6�ac�؅��yn��S������7�V�n#�$Gv��|���s�.Ur�3�9��QUԀm����T�z���z�"��(cN���,�.6�yߧ�+��z��9γ��N����w�T�qZ̊��)�j��Cۡ�̯@���*s q�
f�7"�~=�6�O[��˻�^�{��*������@$l�~[m=�L�/�Z��M��}_	��_��4'o�P^	��`� &��(+Y�6��Mf�D�y?%O�n�ch�_t�@�-�
�%�;_=u�X�%��b�7F����?�ݖ�O�a���F�2D���\k�O��ϕ�k��^��y��{X�x�r�b��|d_�mM�9���G^5H\+���\/7]\�4�f�~ ,��e�3{n&���*���j4�ֹ*i��)�;�Q�c��ۘ緋��_]��C�8W�st����}���A:b-�|i[s��Y�ޟ��B6DL{K�}^Q�.	��r�����+;�;@���=�����4�L�m��D����M���.�Oze�y� c����6격3�)3���z(;�'''�J1<�<����bX!��||�&�[҆&�#h.?7W*�����g�pX��B�w?T�8��rrdI��X�̨������W�+�q�,IO�"�(��������T�_��1��2y?���7撑N;u�:���u�p,r)���)AP~�_f*H'���zUWLw"ڤ�� A�w�; �^��Ҿ�j/�J�z'���r��1���4ei4`_�*O�����LN�?-��ѷ��Iy&Y���#P�� C>c�6��I$����/#�Yȟy/���!���Y����R�|n�B!ϲ���k�0�l��R�9�ِ�{��X�s���m�iJ���̏����Cn5�9�*����)��y��Y���T�FoY0��Ol�A�!����ا���a���>����Ͱ�:\�" ��~����w��=����cYx�Z�1�M�H�6�ߵ6�����c\�.��HF��/���?�{mVz�Yfg�{�z����(�mZr!�y>�(QǼ��L���1+$_O@��p2h�@��.g�CS���{�w�H�!>aT�.<z�'��%Zuq���J;kx"���b�XeH8>���@�5��3ļ�/ۜ+��G��ݻvxw�c���:���阷&'{nfO��t�(e�����n�u֘IQ���y��z ����^�RCuu>_�I����;��[��I�A�5x��y/�ֆa�e�?�����<g�_�R c1u�U<ţ|t~��ɘ#�*,�u>�˗�a�}��s�n3�2tINǅ��!�k�m���M�I����F��-R��с��W�u��D��u���F�������-��xMR.��YUP��>�S&.����o�L� �oW�a�뵬
��0�z��E�m���4��3�xG�ti�|*N�e/5�Iǅ�����6�1���T�����Nh�uq�\b�|���Ad�5t����:b��itd�^�y�3���e�aT�2��B�o��w��.���ר�c3pBd\85��&��U���"�2!q$�� ����u�_�}!$E��`s�~ Yu;����*����g3���lU����x�HY�7���1#q��{�^��Y����חQH)��uV��!�&�6�lZ��M���&��2M����+G����c��H�與fn�Pa��C����u^�_z9�]��Q�W�I�Ǵ�E��>�ң���3&Gh\
�H_o�6;|�_�0�uq��y�%+��O�ڢ38R5�s��jcndM��-l�,zCP6�VF��.���e�`f���p9�Z,����>��vk
�YЍ'�J������f�J�Ϛa��ڑA�7�2�h��K��z__ΐo�e3��xL�h�|�[RRBc�5ӧx��ڕqQ�S==��y����CgO��M�m�H��MB�k�6���s��'�D�L,Dj�e�W�иԠ��9N����~5C_�����7/]�e�0�5:�����I����3��%�_�s��%��pq�z����w
~ʛ�M.*�1d$+�lRvx�Ej�C��U�Ł��^�s� g�&+]��Q����Q�R�%�т�ҭ$6��QB���x�dVG��5����^Wb�ti��oy},����. Kf#C���^��g�č�N�;-���5i���s27G�����y_�^�{���k��߁���eQ;Nz8�S	.R���$ᤍ�Żv�=n�L0��-��;����ׅ��g�!�a��J��^ ����	!v���Yl��0/}HV$i�`��8�y:ZKЅ?�q�!�5����{��� ��:�h]��1�f�������u�[L���9�]0yF�ޛ_��YP�@�-��S�(�&�v��E�3bݖ���~@��nm /�Z�N5 �b}��ثS�3i9�r�}~��ڗ����xjF�V�ϻ��N��SuEmaO���RvP���ݖTS S;,�^�H>heۜ|L�<��~5�(�7�>�G���Ʀ���h���P8Wya���	��I��;���YL@0"�j)\�6�+mn.j,��� ��0{G	��H�����/�EÃ� �l�?�[�k���������4�^)�V�"� Z��L4�����I�̬�s�3���9���d��)��>3fz���"��ȇ���4���&��)b�%�S�yp��%;#Z���V#���k��Z@�Q;'|x�s2qkV`=�ǪU�Q��!-N�7�S)�2&Zk�w��1O�C��#ɻ���=���4k;͏���o9�$�:j;r�N��q��$��'��i*h׻��O��(i(:Ư~~2"��v2�`r�C�~�_FKyܿI\"�y��v�+}&c	�ҋ�>WJ�-���S�#�������
S��9oS��{'�����(5s|0(�S���i���{�K|@H$2_�sz8��ڨ��D:�����w�xٛh;����i����Ww���"���M�ڹO��;��&��;���)U��E�2�Βl�&:z0����z�K��lu-�!�#m�ô�z�#��]�o�Y}]OWS�8��kK��2<9��穹��,8s&�6}TЬ8��W�p����Wk~
�wQ��N=��8o��oI0�g�
Z���E��>�rs���
��P��s��"��=�P6��zZ���c0f52�@5�pJX�@����	Lh�N�Ɍ���-�s�>�8�"P1��������� ��7Mƻ��
�� ?��5<���΅��NY�F��l�MP�̭y��5��y
vx�7Kɂ��s˒�,�?���y�i�Y��b'�Y��>��и
���<��y��{V�w�:ۥ�x8Y�^)�K���dn[��z- D^Jj#g�J���"`1\h|���U�&�U���n�b�c�3��V�K���%�P�mv�ٹ��|�v�tZ�c��HXR���%l�W{Wo��4u#&C�0D0� SL^��/;��-;���E���\%�vĨ���lD������f����6�7�*�q�i������ў��D"q{e���lB� .���3B��nd.�!yNQo+�6�N� �b���ڇʭ�X�Z	@Ri�E�Oz�'m��h��5�2�Eb���sT�I$\����C�_��9���3r�{�Ag�������!JH$>�=�c� ǚ��.�q��EH���K�Ѽ�vv�������s��"c[���E0cx��<=�������-�Yi]�/D��f��S�[����gIjO	0�$��)�+�iî����m�n�U�3C��f�� q]�U��l������S��g[!���كW��5>¦���b��-���U�=O�|��Xy)i�+�st�٦�D[��{�{!���I㠣m��|䳑�Y��sS+!1�z;���c���ov��I�B+��z�~������G��:eu�A�1���/93i�^|��>Y��d����� ����.:�����N�=9�Y�ď��`���m��ϔR�:D?���}
�0�\�r�/��'�x�[�����VK�&�/߃Bo�>`�8�*��0|N����P�4�m~Ox��j���D�M��dKhS%�6��
�O:�K��D��_Q�����A+�:IDHasE(��p5�f�f���8���}�r��)��'����ŕvAn:���"a+>��ig��4,\ml�]�W�J�{�0r�����%������ϟ���á�S�<�5�+�s��٦�H�8��QT�����3��^X%�XE'�r*�B���t�h�7O�e������:�SL��|��d�b�e�������D���#�Y�R��pM�������7F��_ɅDoE��1HT?)l�� �~�l����-̢��Ha`w�IC핡��39k?�tn�Ok|���<�V�O��ҩ���{��qW2$Ș$������0�Ձݒ�,<Tԝa5en/U%�P+9�m��Wdf9zӞ��T�� �ۣ)3�.z.f���cgc0(L�mFy������w��z\�oU�蚹*[&�7Җd�v�,/� 	��M���%��^ p|u��a����Bj���9$�]ԤQ�9iS�.�M��H%�}�p<S�rᑝ�\��G����9�%�E��%nխ� c68� ��n�����N��&���$o���U�C��ڣ�/¨���*"�W�ߴ�J��]�6��쾛�}�&�$�*�Ϲ�yk45�f����lx&qv�
)��%~��zG�h���H�G�ܢQ�9ܡYq��޳i��N�g�րm��Ja_���V,��.ز�6P@���7=���T��^��ɾ��런�ݝ�.��:G럏��
��*ͯ?�f۔����z������ŞLz�*�sP�Z�ZD��*����+���S�!�n�HIoFZ�}%��t����w �x֒�r�/��3Q���݈��l��ɠ�'p�'��a#/���x�x#m1�ZHz�����k�7y��w���Pk��ů���Zo�S4O�����(����b���o�R�vTq�"�d=�;��Mu�.5,T����O?Z��i٩_fǗ)h3���A����J�d��������F���B6	���PH���֌)�q����%C����?s
V%<M	�R�4M�	(�L�2R�W�E8����Np��>�6�|ʖ�b�W��P�$�nb���bVD?�5����W�<�#��N�G�҂���R�=�VFF��A�{!>�V��	�x�3Pϴ�zv?�z����l��bY�e��e���3r��@��*��]ϤM��w>�Ƃ]��NSS�5;y������G9W�G]�ȸ��=����(KWAA��Ӆ�;�iaq,�@�rL#�7yS�|�����۹�� �!����M�����$;��Ë�E���Lo�������_�f�av~�[w��4.���4��U��,Z���'r"�"�څ�8�d/���+y�ȩ6a�l�|�<b���a���+?��Tv���p�W�1�2b������.�li��6,�󋜄LU��@g�Kk�=���h�]z4�}&3�� A�FC�.�"�oV�aȽ�#�,�ܽ}j����]h�E�>�(��>��J뜜[{�L| �c��>@=CV̹��Lc��|6���_�c����I���lǧ�u�2g���b4�"�Ԙ<�1>���a
���cC@�d���XL�GO�7�+2Wg�%�n��c� �Ii�dN�.B�F�_5EO�L)- �9Ae�LP�W~k<Rd��PU��:���	�W�[&���
���'�x�?Ak~�������A�7~"ծI@!�V�s��@�9��y�s־���ҫ������;��� ��Q�V
[��8/A�5o>M�V6�2�bڐ]���x	��n������O���ގ>���Z����M����T2H�|�ۑv��L�8���i�y������ylz$`:���	D��/�mя\k��~6Y&�A��c�}&!jQ�r,�뙴�H��rز�V�����h[�N���	?�_���Q��EȑH��Ǥ�p	�Z�4��A��>�tc9R�g��맛����*��n{:�-���*�?,������� 8����<Y룢���(���"i�5nQ�7��)�n�2���>]�@�O�\������Ԃ�����踳><�ʴ6�JUԗ-.�)v�`/'�[���'w�&��fd��~�<�^]6��4;|��^fJ�>���Y�')�33�����b���<)�U���~ŷ9Q��93ɗ�y+��+6�_��̾�1Q��6~��_]����U��2�m:C<���r�|8h�*��0�7�%0���w��(���0���Ű*���{ &\'��Z3�����ui��+��!]�&R�E먀�ϸbg����ՉpK���*����@���ŀj������I����.�#�����,�ǯl�=��϶��zc��B6��0	X��;��o��yt�i�;����b\h(:�I���>�K�Up����[��n�LJBY�?kq@������|�On[����A��"��,�-1J2%;*&�0�rY!_rs>�.hG��Ӄh�w�Y��.����vo���3j#XM�x����12�/�oX=�Q5�ߙfO�'�@tk���}�)r��#�铟u�{Jm�0�����l�v&��q%@j�/�˚��*�mL��Zu��E|y�Q�9�(	�Se�tK�~-.y��&s��kf�5���Ռ�'�uJA_�\�����˺��O�9C�Rs�*��|��qئm)h�on��h0�zz�y�d��\w�sl���}7?��F��� �r�H�ix/�rd0D��=/�\�Z?�!h����v(2xL0�з��H��~E�~����p�NiΫ��2�����%Y�ۚm���^�&<�C�ACC�������/��N��Ϗ:d�$�nI�5�_��[�������!011�k,�gAfI���+L�i44������@2ᓍ'�O�Gjk��G�Jn�u��|�q�Glb��b���)�7ɥh��W�=�f`�:;+����37/�t�M�{���XK�M��H��[�7W��Wi"�m��[�A�X����WI,���O�H����6������;���⃚$A���?=
Ꝯ��\0?w�Rڄ��~�ԉBƑ��wXE�J�{_ס������N��y���6J�E�`a4>Ʒ�e��?:�)�҄�� �R'�4�g:�TA9�|*�^ �r��Ls���zK�j��	 ))���3�g��^�(Aw�L���؟R�۶ʵh�l�+Y����H�T"���Ѽ�� �Js{�\�#ONN�Y0l��qԵ��ǭo���Z2�AR�,e�ǮH'��T5����������م�X�Y������Ϙ��s]�WX�W�pc7t�>���N�"�׫u��X�h����/���G�E0�K�骈��;Y��c�T�Nn߼uk��S_��<ޓ����n0``��|idC�i�Ѵ.�?��9�̷c\\_e���e*�������*�P�ޤ���}O1�Â9�����%�y����»��@s��J)H3�({]�r�qBD;��Y/e91
>�Կ�n���q�|ً������&�_�8E�ggh0�u�߭��
�R�+q^��E���w��L��p*n��+�<]��!×�&��B}�����M\�Aں/2c�f�m!Wl��Ni1�>���c�vT�z�o\*'��Os�(�����IK�8Xl=�h�\�Q��β�W��]��+��![�Y�W�D���4].��R�]����U���l�V��=va�GT��&�	��C���T�]���kpaƠ�-�U�V������B�υST�&	T��O�O�L��"@`�s�fx��F�l��U�
i�4IJyi&*n*�D������M��FKV��μk�Y�,u���33,�)آ�'<"�¨~�c���T ���M��V��'�?y���g��-�h�!e�^����SƏy�8b�������;z��D�oF5{�<v݁���fˢ�w��=��;���X���?4Uh�N"���{�Uvzf�[G�sR��Z����Q�,���B?��D~�iJ7�mɥ�x�ѯCt���ă��re�Ptu�b���)�ǅ�~���SƁ�:MQ���������젡�z�Pp�tt�|rڟ�m��\�Y����wл:_��:)��xF��!����Nx�g>BN,{��C�л�L���J�0��)�H��	�[՞��~��4�١�9T��Q^[�d�Y��j|�|8��n�� ��E �?G��<7,b��c܄dM�gLOw��u���ӆ��ג�f	���Gj��g��һ��Ţ�]�(��]���5��TQ���F'�caC< �΄@+�{�I97��H��ޠ�>k�ڠ�56g���XN&�^��ˁ���Q��x���rR0{���Ѥـ{ò=��>b#�@-ǆ	�z ��K��=��\���������:�(�,۠�������'aE���ܼ�:���]dß�� �k���'b�/�x\@���
�֬ճ�������,��O%8X�	�z�����W��&Y1��Y�����î�H+�����^�8���]wQ���;�(��/��4{<�Z�J൙5���H�]]HQD+��1�T缷ک����!��g,0wW�T��v��o^�ރ�v8?�0��5O���`��������z'���1k6)|��-����������i��I��2"{�5�V�_�ޫ�bYȨ7���6�M�2��m�l���<�pRٯ�-�f�#�D����@����k%{�\K��n�N��7����힥IjR1�}�6�at�j��V�����P��N��`w��t���P�ʿ�Ʌ����n�f�B�����bg�O���_�J�t%��[���R���x�ػ�q�����}_tM.��jh2K���ėe���}6��xp��L�q7�xЭ�f�x�#����&`oD�ۚ���Y]n�F�&1Sā_Z:��`���Y!���n�ǭ!�Y��'����Jׇ�R��Ҽ��ge���f7L"�.u���$������}������I��m�k��� ś��)v�����A��!� Tmɕ��ə�����+��,ꏓ�����%e}e�zo)�������Juvg py(����+�QVsS�d@`�g��io"i#��}(�XPk�;�U"t{��R���W_m(�ݽ����v�eх'm�b� t��qҜ�k�N(�K�t �`��=|�@~����J%ʁl+�Wj%�+�(�~��<o�6s��Nˑ�3 ��t��~�S	_-Z`ɻ��"��Y|ڄ���#�=���-���@����C�C�9�����2�qsȟh���o̾G�H׽V�n�� �5����V��H9..ߎ.����@�)z�?z��`5���ɡ��z麟#�$9�7��dJ���쓊���S�n�	�\H����D���Q��9�6L�jR�ν0o���s�es�8���{�7�Ǽ-H�"�@����c2ls�q��<���̣�C�y֚�.�Z� w��~�:V�iB�k�+�ř	��u����wq_�_��ij�R��d��6�_�q���b`W轿�Wb��}ŧ|��hm���H~QY4��Q��҄p?|�����W��m��<@�+�>v%_99�Z��uҘ�+2g�B�ā֨7x������p[s���2msю�,}����dQ�{��Z�`�E��Ϗ<���T�`����s�wR/Zeھ��1���]D�5D����=��B�(-���[��Y��=�����Gr����;Y��K,_9�C��[q��PQ��ܶɐZ0��q_޳�1�$����󛃡~�	����
�J"%���9D,G��Jǃo�?8hIHb��0�ha�s�&}?���}�n��Qz4�����G�]�X�*��@:�9���]��ځ�����iv���'�j����'���1P�d����	�K�+AUI��7�����}�t��5'0�r�%��7�'���M��5�^�8�l!���5,@?���������޲��f���f"4m��nŮ��VZ�
�R��K�uI��Q�bd�I��ݻٜ,�F�3�\��e��0x[L
����l@+�M'@%�����Sg��6X�Y41��'���h��s�O�����pL�@B+�\� ��z������ۍ4ȥ���������%ϴE�5{�'֯:��Ka�^0Y���/_&�a�n���aެc�~X� ���ʗV8!���R|o�״_+�.�7!�a�w���P��b�_B�*COK֬-��5��y�K�@ɑ�/L SEoJsY?��'B�r|ʔ�MB����՛%�?�<R��[Y��)���!+B�tk�2\)���~�1�r�����G���&_��[�7�n��]���
���%��s1b��A:е{�J���'��#���0�6>���#+Õ��Y��e^�AiZ)i��Q�A7�wTbc#ˁ�),ݭ^��6��@������jm�(!-=}_S�b��Y�����ϧyS�e�x#Ekང��Ox�X�繿���=uD��-��d�o�Zg/�Ĕ��Mu���mut�����e�潆�l*� ���N��ȵV�4<�����7i����b�$?u�i����c���Ƨ(���,x�6Yi*ΨL��Nȿ���%���b��rt�/��v�I}��b��fM��1Dv��J�~^����U8c�KtR�Nq޾���&8/Wu��W�~�/Q,I
�O�M�(ǎ��>�I����?=���h>�E�'ᩡ+"\����c�Բ����[�����U�՞����w�_���H��I�8�X�E_�r����eܟ@5���EÚ���w�>trAt&&&TTT�ד<����;'/eo����clp� �����U|��r�^�`�bo/���r��
����fX�{��B�Eg�\��QRQK�^�Q%����(A�[���v`߬ѓ�}�/�:�Z�M'�\�jX�-ʺ1׉Z�aP�	I������dZ�_�bēy�P�&����+o͓��`���2`�����*�jy�@/#��*����	���_���Fq��)72$�(����L��$h�h���*�}!.Z��4;�� g�tz���/=��b�ł��n(r��H��bC��i�k{�����xؗ$��Ό�����Zz1[RR�/�Ӊ����N��j<w?�76�����m}O�(iM�$c�4lv��xa:99]��u�nmm��T�Z�w������PL�	�ϕq�5gI�_7���m�}���ƴW���e��ܕ=��K���c����Cw�,�aq| ߧ�`���2�y��+��i�䜈t��t���t�&�� �~ɱ�Lw���I�'�(q�{-0�Ν�d����oWI��B��p��w�6GֆB~�<9�Ώ�C!�X��o�DҢ4��B�s������X�wAHC��{�v���+t�>��,Új���r&uglܺw']���G����\}��ި=!�&/� D>A���ߧJi�*U�a���/�8�D�ar�ÿA	_��K�<ل�P���K��
X�yNN������l�靏�+U�t���U]w���\�^*o�¿a��/z0�'8�Z%Қ-�%��y��2�߽�]-�ekC��Ȣ��ȗ��!�!$97���gg�H�e5E
_��tϵ�~���]f�-R������`��O7��e�ɥ�4�T���9�ס<�����Ofv���e>�fs���>�5�10o!��{��\1I�&ݸ�a�3�3����3M�I�������y}��*���4x��h��bg�5��y���!�鋼�P�����1*��ôP�z2Cզ�JԦ��$~l�䉳�k��z��s�M5P`9�����;���U��n,+��w��k?'%�����e�6��5�eS����i}�;���������-��B�@�-:�***��I�P�I�2�<�28��r�>F��M]�w.��k��Ƥ���+�'�T�Dh��l����UT�s��.�z�i�b�ҕZ�����9�;�:��\�N_|5>�AV�Qύ�?�{\�q�o��f��UD@bY�-͟v4=re�U��p����?��c-n`���A�[�/�7�l����DԮ��KJW�A�U����L�� =��U�����/�Uf�M�$�q���'�X�;!��u�.}���;g�.����Aŷ�:{�N�L�7�1�=�4�*��h��m�x7�,IÚ���7x��(_��O0�=;�xѴ���#��m���LV��Օ�_f�؇���o�!l�3�ey����ϴ<6��p�[�G����=������dct���%�vҩ]ME~�l�x��d&"H��6��f/�\�0O��"H�r��(����oN���qa;�Fe3�����فi3zΨS�Cam�c�[o;#�$)�;oK���{�rk� �E��B�_��.]%#�Ր����op�b������w���`F�XUz,d�d=Y�MA��U9,Y��
�i*����[��
?nE٣����l�&
Hgt�X���dzr?���YT�}5��$�,�jK�q� �X�0����9�յ
ʊ﵍�z��#,8������[�}A��M2��Rx������a����h��8�����t4+(-�N�q�TkQ6���t'I�(��V��u�o�۟@����	�����1���%IIII�38Jc:����6?��}������S��=�$��}���>% ��|{a��OK�ge�
�!ڃ��Q�:�pw�(��+�����6��6"�)��(�/��;�ے��urPn����D��)�Dn�����b��z��B�Sb�VDe2?u~�+���J����!����$\"\�Q���ř�ր^��j�B����Ʈ���ꃜb<�ޠ���XK�}E���Jc?�cW�}�$��#E�=��]ߛ�n��K�MK�"�	��nO�E6E�'���
���h�Oag��s��穤T�>�y�ƒ��JCkJH>�����$䭇�"��Ի��Yn�>�.�r�/8�V'
����;����3��[�t���w&F��[�?�/��e�öb.�ޤ�[��>�[�-�
� ���I��.���	M�,B-6_^o���L�#���kЙ$!#9oiE}��'.��-��g�$* P���m�z��  ���/�!~���ET��M�:������F�� �ae�@B�ٻn�/�Zo�ԏ����cL�M��Z�;M��P�/;LS�@�F�*q&N۫��S��s�߄��b�M�6��7�\_mG��?}���.ķ<��̌;b{�c|"E���%���1��	?w��k3���@:��}��v��[ca���rK���1Vq�3R�D3V!��y|8v_��q�pm(R��;�!'��_i�h�`Ӊ��u��6��!p���VVB|�
e�v"�\�Pw��>Q_U�4ɖ�����4#�����ᓖq��
&8��Y��4Uz�p	^�����U��*<�u�᜚e;t����C����
�����j�$�~�F��T*�+Z�֮�J��ܷ�N�o� N�ԏ��eY^�]�Ԛ~�ؘR���`ȜS5�/����FXklf�S�������Ӏ��Ml�/�Ы��>=��oMT��l����r�s6�Hh�(Y_�թ����"�?�5�h]m�?���\�Z����o�Ŗ�����*�lU���ϐ�W������,��� ��4��.7��)�)�1/�ƠUtQ�
����C*�#���=%�K�P�'G�,��/a�M�Y ����lj�~�l9&�l��MV��&5:�N�ѡ=_�}$��Nﴣ1���_��7��Y�F�x���|O�J��:�k;�R���������`;����66���>���`7˝O(^{��<�ۓ�����U�௓��*�B�^�q��9�����N����I73��u ��s���|"���NM�c�ۨN����/~�P����f6��ÛR�LC��A�Y��*����G�A�s�f�����e�G�䌱�h:�?����9�5c���5g���%�W_$d��N$c#2��h�
�DX\���;�>�rĚ>A��Uq����:���
�頝|� J����Paf�����'���*�*��c �ٜ�	�`>���f�F��憟Љ�����g��·J�����@��瞥�l���Y��dț�D�;�d	ݼ{���� ����o\��4^[�S���?Try--�4>�����ƵFAmm���{F�?��F�vvw˼2a/3eھ���'��.­?$�Ey�r��±�x2�_�;�]��Ѝ�/L�h�~��[�����f�z�>f0:ϩ��L�]���my^�a�s�,vg��}=�"±���A)&����#�jP���uv���Ez�p�Y���'��:[s/���.=�p�E��=
�q SRhQp38�3�I�͑SZ�q���%�9�h�Xô4�'��up*^�R=��"��r҄P��^W��h{�e/�F�b���Ks��*�o#�HRE�s{o7N=��~ؖ���I��	���‛-��������8QkzN��٭	��d6tz^v&�`ܹ��e~p@�X[1gX׿= �����ޞ���?����oq^�%f���V�լ�W�߿������]���������S���1��Qm���8�)�R�w
����wEw/�)��]�C�νg�/��/�w��=��y�0��1Z���u,������a3X�����:٨��O�^k��솒��y�����<�>���&�d�A�m�C5�nOş������J��T�B��CP�_-f�CvZ��'Ũ���I.[|P�Ķ1v�����d��#�#bC<� ��t�	ۓ*�<^�Z���M�ԌZ�����g�$檌'{����{�`�����D��,�k�?�F]M�eFw�.d'DC�I����@O?̠RG:+�T�
)���h��|�w9��}����h��u�umr����>�CJP��J[F���[}����Vp~��l�{��ٶ-�����]�!��Z�������_Ҧ5����/f�m|÷�u�� ��Q����A χzs�|��z�*�O�ը��,7R�����D�[М�`���\^�D�Ed�Zzѭ|����/}�����������i�8X,��>t٪Ǘ����4��%���m���	���Ĉ�]�8�$6G:xLXn�xPE[�J���b����Y�|2����Ss�Z#6���ݩ$�+ڕ%LW j]�0k���S�~-{����'f8�mE�f;UDw;�:�[��F��`3�N_$\3�@���Jwu����2��y0dc���p?�����,//�Ɗ��2��Ӂ?��l��5�[�뿔u���]f�T�, �OA��>���v�d��&@w��O1�C������WU�w2wJ�Jc�gTy�<gưEf��g���%��=T1�{ԑN��\,�9��B6r�Ǟ���q��ݷ�5�_���(1�V��W<E��ր�k8!c-a�h�	�oa��0R�nK��=�%>�M�w�f�lV��S�Y�]9�f�#�`����{�ScW��(��+֗vq'���у_c�\@^����h��"]2:16���
�F.�'1yr�HZ��;:�^��VOT-!O��JY�{��\�Q-XB��/6���	9�����m��[�6����<?Y����r���-m��Ym;.#����Ûy��f�|rjJ��C3���F��;<?�I&}1���)|ZT�	����X&����VA��=#b�W#�Q�;D�4�k�ċO�R�P䲼�:�6::�ҙ���`�&��bm�ɇ���VvW��v�7�Lȴ^´+��f�ؾ��C��]���G3�"��n�Z_�>�uu~�: �M�$�o�=ɆP-�ʙ�C��j�Q�C�Y��5;0��6�� �h�ƈƇ���xH
�t�����D��� �.1s�H/ �\~ρ�L�03KGܵō��xiGƦ3kU(��w�#wf�s�u}��\�)Z_$0ͬ�Ӿ��\"a�8�����mxv�̿�b���x�ҍ�Ņ�������k+���^��Uo��7�9��_E� ��`�������/��8;c#�>i�ֽAt��^�U�E���i����l	��6��=#Fsd$>�RS,�_I��gV��h��m͢]�G,1���z�!���l����lܮ���9�3�~��fn���z|�����&I��X�F��^3�Q�.��I���N�|R�c9=�i����V',�@� ����PG������n��g@��y�K��u�����8��z;3g3�����-�\��0����׹�k�;":��cv���b�D�Dp��(;-D�
l��]�0��ҰG��9�S��xƌ���r�ۭ&V )�c� ?)��U󲽜�IEbO�*���6v��������7_���������J�}��{��Q$<�2~�

�kO��зv�r�� �]���/A�Zo���{U<w2����=���E�@������%�Yh�����z�����B�x0�3�J'���:&~�ݥ؎c�������+�@z�p��f�Pn/��l���%fr��	����l��}���0;q���Ϛ4�e�Cx���Lc�LB4C5��c1Dv-�5��j#R2~�m���ɡ����?�;�4ֿ$�k��O�h��s�Y�����:Z�}���'�uGO��>��x���jmsh-G�]#��uz�+v����sO��ylw�ܨ���u=X�v{�5�B����H�������|qc;��?���tg=-dm����� �WPzŞ�{+[۾��o�K��U���	�"�*	�B�w�xb�����Ȱ�ȭb�Ö\q1'����b��9���Kو��XTn�@	�]n�w�L�;�Yg��q��1-&���ӗ���]��p^�S��kw�Bn�u:��\����F��]&Jt���׷���qWVr��ul$�u�d%��sI����Qb~kw㘗�Q�:��L�'�Pg�=��i@Z2�v�O�����ǏbL��	��m����w1SM�A�����G�ߩ�Z{|j	�p��"pm�|�}t���I��G3x}�C�V�T��QV�Ħ&��NX����
���������WB?|낕̎�E�J�v�Ը�M�3G�̓r���,}�j̽�a�Y+������uFGGk������wܶ�n<ݮ�93��l������]��f���kLGGw>�r'����v��#�/����:"7�K6g3�(l�6��s���OZQS�"*H/�c�Rk�nP�|�1�XK�-|Z�O�� �9X�Er�i/.����m`�~����7�|��y�el�I!�����A��웋�2�����cy�-�r(�o6��8a�Zқ��՚�M��ԛ#����Kc�},L�bs�ab�y8D��ƕ�r��%��r#���>�L���ݩ���gPt���s#��gvBpi�t��r,\z?����K�}�ݎ��Tk�DgH�ߠ
�2���ʫ�fbN�½����P���Ԯ���������mB���v���e2|��`���s�*���ƞZ���)`_�j��A�J=�Hʱ��&��ˣz��ëX����WNN�k�f=�%���B�=�`����k�����:�?����1~������쏡x����ZL+�-F䙗�c�=:��d��d)��^��sdt�Y���Q��]����ٲ�ak^O��G�Tp�PP;6���o>��@PB��C~��=���U>[C4��p-�+Щ���kl��|��$���~g�%��~�d�T�#��1hD����)�t�s��m@��*IY�9���\����cF��jS�7�]F^�tur��b��KS/����~b���c<�b���)2?ÿ�5�`0�M���zYR<H施6}���*�9>��ǲ���(v<��"�P�S�润k��C!�v�����FJv*2�"�R�^Tajcm��S�+l�U��}�/.z�jQ�#�_�M�+S��b�]�߰y����y�8���6ⵇ�hq��Nq{�tJ�>˗o���U+�e7��/2׷ �)d
�^W>�e���+ͼ�玦�l��S���<h��⯬���B7By�n���K�!]/�NV���t������@
T�frIgl�3�����>�Y3���!*&�Y��[���?��cf]�06�����9u�pf������� �Z�ԃ�^�Y8���1K
e>A����Lx&!�7�b5�E��KGh^.�ƍp<�{7յ�@+)�6tϲZ�=��h��"B�Y������qoX��WOk��щ ��!A�=D.X/����¬����3��!��z�Dwr��+w%��rqg�`�������-8��oQ��ɤἝ�>�`W4A���e��x�q��S�O�MT�LA�iY�� ji������Zy9���:%�Z�f+���w���������u�DSItEm��$���j��6����
$�rk
d�6�N{f˵'gg�\���1��8/)�/�V�W�%F6~�\X����rN�-]���b	褗��A�Tb�}PEM�]��A����g`X�Y5<�nCC�&���A�C�WA��V}?�z���%H�m��%$"���X��U����\A���|Ꜯ#B̒v�|Wzʠ޳�e��^S�� t�#�U��٧9R[��[��0D6�e�>d&��a�ha|�x\X�x��n��sb,��7��ǆs>;�U����)���+fC`\��V��B③a+~��=J<;�����p�u�6�F����E�>�����6�d-��� �α}���˴��4{	��y�)�)���IݼQ��B�l���ej��w��.M�6��ZS�΃n7AK��[Tv�@��2����ȶx\�|kp��tC�>x�6��Lɻ�kΨ�=�]"���v���"�5�
��#�T֤�5��HuW�ˆp�(����J��������B#`Ygҿ�y6,q����r=�j��M�b���w\F��ǋb1\�/V.:[vE��3.�*��*Cqy�F/�m""Y�����MY�����
�f�!
�y�Xu��,��ˋ>�V�o��z�=�	9~H������a�h��$Ѣ��p]�k�|�6��v���}ؒ��?a��J�`8x�c>L(���Ɯ�.
��9ݹ|���S=���5wM�U�5���PY���ExV(��/=����~�m�n1�$h/��0���I�c����B�c����.�ZZ���1'T~�3�*�5��V/�u�>fp��K��) �a�m��a�ƙ�&ۛ�68�a�`�ה��M����� �E�*`PC�ɒZh~���;)���`mԥ���H�\���qn%��4�>��y��S ��t�<
r��=�Bba9�?s�t�)����EO�0+>�F+�����n�����|�u��4��3a�௥�q>�1��c����Iݦ�>����F렙���lF�nn�F@�^�)v(
���T1��sv����i�����2=QGG�(�ޜ`ͯ�bg8�D //?_m���}!�|y�?=��薎[_���;������Ӓ8�m�8��!2!�d=f|T[s��VR?k�eӓ[1:��'�i�xqs�8��(8��7�\����F�\���L!iNO�=�s���VH�s�2��~�U�������(,�8:�݂�z�SO�s@a�����/b�e��~��tˣ��mi�i�K� ���,h��r�4���CTe���W���1�ќ���-:���4|�#��㳌�zZ��ŀ��#�0�_�dG�j�?EݼR��ѓ�����y�b�ع�"�h0�L�b����a|2Sr��|:y���>��������`��*����1�_�0Q�w����tކ���_g����P�ڱ�1e�X�&z�r����X��MS�]g�nW�曝�1W���� ��j��w�_��.�-###WۭuX���L����wd�d)��q�WZ���/���n!%ǣ�77��k���'����Sē@!���1��'j��j���+a`��;j�瞾�P��q�6����"��Q���r�Iq<K^��0uw��n ��
>1�Y�NvY1�R"�,�Y��zu�@S'3��
�/ܼ:�x�~V��J��[ƞR?�$[3�1|�@��Q}�{�Q��;M����V-�iq�����ؑ<mU�, �DHxcܻ�I���ϕ��ޗ?�Tvo�k�Q7O𡒟WO&7F�\�A�̳*4�j�ko�a���2�\��ۯy�b���t$h���Z3�=�sV1�x���f�x*i�[E\�ϲ�M@�;�CW��Ӻ��z���B� KΣ���_�Ɇi�P�I�o%�;pR?�]�5R�^z�uT��Bjj��k>�2���O��d7_�� Uo�$��Ap�
��	�\�v���Ԋ�Z���X��[�r����imKM�W�rMBY
����L��}�8��QX�U+�v��=j~��C�!68�ĸ�������vY§��^�������)���/>v�A2W(�,����>�tA�iv_����AxR�U&opL?;�p��M�5!K-_�Dk�8]����zr�b��G]�<�r�6��19.���~��q $c��FOE��peQa���iC�`[��N�>��}���n|��A�F�,\��of�����ӆWU������G��	�,�f�k��[���n����-���(E����
S^�-�
9�����B.��f��������Ɉ-�Y2]^T�rvd9^9�D�1�}�v�#\��;�$V�>;����j;���I�^�O=�� ��cc
�WE"���_hj�}��Jk��t�k�q���C���wGR$�6��?v\�n䄒�)**��\�	�2� �4�i��!/�ȿ?�Ujc�j2#�������Q�_�hj��W��'1T�d�;����A����y��y�PS]Y�\ۑ����+zk�+��+����R��|C����Ib���~�����(�Bw�Xyj�BTհ��ş�D����͒/B�!�E�C=��^q@��J�Œ?'��VYқjxEQa�F��7?J*��_%�ɉԆ��y�z#o�-������7���(��a�`��g���Rz+��W����l}5����u���0�E��{e{sȋ733I�),��e�kb1����A�U�����/�}�����@%�>%�c^6�bT������b��>�Vi��%���hRx"Щ
�Z�����q�}�x��)��v Y���I>���'d��S�X�pg(�8��u����~^�n�)33���?�6���rr�5~X"�U����K/;�7=�HX:|Q�(���U���qBN�:���w�+�RdWX�3?��'�Z���ua�?� X����Q�7=
.�hP�tH��E��nK|��� �H�
Y�Kq�&y�����^y���~����ѫ��A�A������
?<>(���m�c3)������
�'NzPMa)"¢���n$m9�/¯����}cm��4h���G���[�r!��~nN�[�a�͡cS��g��;��I!AZ��W�w�6B�950;��\��;�=ŝ۱r�z��~����y�xo���)�ԆQW�7X��N5�%t��HZBlؕu�+��\�<e�!��VY<8�{�+�5��ܙh�q�x���K^��Am��F(E_W�h��^���&�@����ci_�s�I����/��F,燅3͛{zɮf_��x����a�2 ��T�$8\�R's+�;;K�^���	l%�-> �U�;�j���0PxU��p�(Ѱ����7u��$�k���k�R���}�bB�L��������O&�sx%����R�^�b�#��(��x�{L�k����/�>�BN�[��w�z�'kvWB�+x���Бm&�z�L�,���<�hI#����ŋ��c9���
Z��c'V���oS�93b� �B�ho�hٵ2�4+`"�<%�V��B��P�M�C^��B�{��6�ЦE9<��X*���/v> ���A�3�|�YKm!�J�
y�o0�'�95=`�����}n��PL�d����/���2�'ÒN��sٻ�bn~�p�5o�ג8z�\��� �EQ!U��Q��K��]F��O����f����3��G�	����� [y��g�_?/��xu���x�wJ�R�z�?I�)���UhRps,e�Rc�S��)1u�8Bmĸ�ټ����Ä�&m�nOs�&R9�C�hQ�&�>a��v���_M���ry��{��.x`iw��ls�w��W�|���ؙT���{.p4�.�[�����s�'c�����Ly�'�8�{]=tT�b5�k��l�n��)��G�xŴ��a���8k6�]���cz]�o�h)���v�Dz[oTVD�j��5Q(�-8�o�ں$��)Eˢ�턎������&\@�Gqa�/a*�N�#Z8��c��]���ʩ��Nz&���)���K�.�z������� �����1�RQQA�+��1*�����gR����A���;����ۭ~�g��a���3��{p��B��+�y#���BK/Y��ͥQ��p��"{���!5��0�2�4|4$,�-�Mâp�|Sp���(�Y2�>Uk��P��]�ݝ�%�_I�qL�c����R�w-�2��?0��o����W'*J�Z��cM`�H�(�
>otlm�V���[$�$uM��T*���ě��$�՚���n�����[1b��F��&c���d���oȄf�7��ʦ�x�;:�EI��ѓ�j�Ӽ&e#�7}�<���wg�Wh���;k%�ύٝ�=vw��3K�h�k�81<r��0�\('�Gɻ�Ab��Ko�3a�9�r�P;Iu�9�BT���#j�V;��B�S"�k��uL�}&O��~�?��s�&_o�5��m$�&��hr��v���b�8pMu5�+����|<���?�JD���75e�ե7��y/95�ʙ����ֻ<���}��в���bC�_՟��g�\���#�o�&&9rKgHj�qo#Ҡ;`��c�0��Z�T�����D���,"��ē��>�g+���n�	��QՇ���BDwS�R��p�H�> �����v#�{����[/ªKO��<&ˢ��:��p*Vy�k]V�~��Q�`��3�U&M����j�0�v��9��$b�8q�`��X2�6lL��FsU_t�Z�R[U�g�8�Q�	0PQ����P=~kR�[���+#�N���OY_�z�f�=WQ���6ml<K���ey�����K����D:Y���è+><O��h��~W��%����>f3���\���k7�4T����>����a�E�ٱ,���gB������.�-��]��X���'%��I,������q��c�|���{�$�7\o���]�j��ɤO�� �4:�ǆ_��.�=�%O`Y[Qs�J��J���攕����AB�L0�
H��Mа�4�T�G�W��С!EcK�,<� ������N�y���oZF��9��IRqµ���c$A�E����^Bg��b�U|�ZpNI���}�Ksr��j�P���5gn"����_s�Y���}Q��1��D&�gm�gjI�}���ؕA�zsE�Xѕ_`N����8m2�g$?@w%��X��Mvdg=�w�lKQg�� ��%9��C?7_���I��-qJ�C�Xj�~;'O��/�W�n�O��l�5�C��D=dEA�k�l�v�����E�B{���H�\�?~�*���"���n^�Nb����6���.����z��+���5h�o�����W=ł�JD�ՎGdff��lQ�>P���'t����B_SJrKE0��}Q%��^^�T�5�5u�W�UrC�������p̢0>슏|Hߏ��^�����q���Ý���Xn �݂��%��ZF.���.�=�wR��[�<k�^Y��=��[���^k��ph�2�{[�8Wo�q�K��fl��P9�Ԩ<S����U]ƫV���@��!�8�ĘE<d��w(s|�/�;x�d���n��U٦>�T!���R�lƁ�q_V�l/��qTB���O6�ؽ��L�nU�^p�?�u��	�LZ�\n��P���yY����J�9��$#[N{�i���<�� uE�$�PeL��ӆ�}"򞅤�.9�g�ڸ��Y7�$\��n��g'��yB����B�b=�0Wa%3���	E{�b����_#�[1"�G"0&����s�,�c�g�	/C��X���&���y�&�D�{�V�_�2{��_�VlR���}3�C�P�s+�za�6�	�G{��V7]:^�4��#Å��D��{5� �ʄ'T_bHqB�����h��#.k��JY�����������������?|ĢT�q�Y�Y��{�Y�̬�T�.����*�g'#�Ã�`)ʳ�9�P&hw�%�����}�L6�w��]�ID����Ҡ���ZVғ�*�/��r�ݞ�s��T��E��#��;L�4p����50k�إ������!C�dQ^�a�?� ��S��f��6xX��$�sz���ɭ��)9H���>&�fTK��h޼$K����;27�m?���s�Jִ�d3�`��E�W@&�^�A�8;b��$�I�������~��Fxµ�_��c�;��8*O�K������Я"�p��UH�=~�l�U���K5!�q�>S�v���jpN�I���,ڊ��]�՜l�n<�ϻ�Ӎj(=�9]�p)l)���\i"��Տ��-�H��w��`���ZgC�_:X��Cu��L��!^"4џ�/U�Ju3��˵�Zwq6�c׌��?���,n�3Q:!��t�)<?#鷥W{Z��+9@���M���<���_ް�?5��i~_�W̏�?����q���H��8�n�k��(+8�
�V!<�ŵv��3{�$�+���ր�v}���$�x��]�����1��J%��>�HL �լ�^�0�E:]����Vp�--X�����4=�,�?��֮�y��{��~;S�K�N��`��ER��wz�(Bcm�O��D�]��]�ZJ�8[�������4y �sq�M���|��Ō���o����(�b����L_�H��{Pn�~�W|Q���.;�B���"�E<���4�=��w2e�*@�`�0�'{�!�3�t��ki/�'z�N���?�)���&|d��A���ܾ�L��8%Q0ti����5�5N3'r� �Lf�Q�`������L����R�_��$���y�E�����?Ʉ���\�J��O���"�Eíp�ȵ;b�|�U�	t�Շ�hw�!ֆ�׶�o㥗�B#� �p*ڌ��{����)�Q�{1Pu����R���9I��q=�g�3��4C�ckVh�2����2���C�i]�����?rn�|�3a޸����͕e�e�	lcdg���i9b��f:���I!SP����~�ӞB�vc�kYz+k+���z�>>>����@!���xe���4B;D�"6T�E�N�U2���U��C��<�{e�l֩J�h|v��g�L�~E겿���>>$�T�)��y��u�l[�<��f����^�"�~���]��:N8�3��r�_�^E0�v����d����ѣyHVh���e�8I�b|tkݨY��j���gϪ��*R��0�"]t�;G�E�#�>U<��|c���;77��{�L���(��7�,�]�Jf�?7�;�M	��w�;BGr�3m��1v�.ܽyL��9k>ܠ�(����O1����f����]�d�C�xg��� ��扠ѕҪV7�����Z��'�����5� �i�~��/�������v�	�+7�T~��&G(z�YJ���"���y�嘀�Sl-x�c��T��l����&>ׇ`�t���n`���eZȎ~������ D�ү s5���L9y��8���5�̔E��߃��+9�Zo$2Ђ�%��u�$���
�3�ӟ�����ۡ��d��VRD-)8Ṵ[F�᢭��ߏ�
�k������v�,��L1����:�z2���5Va�f�8lF�J1	����d�[��MSq
�y�z6�x؆��*�{�_6�}���Ղܡd<�u	[.@�;���c��x���ƍ�dY�|�������)���ћ�Z���-)��,7�#*j��j�d��8ݢ��g9MD�[�mK�VO�� 3�ls�~hx�o���I��m٩Vț	<x���q-��2p�$��!��W���B2�cO��������?���j��&�}�a�:���f"nkg���*�'3�/�E�t���I���p���̀�����~vv*�Y;����|l������	!ږ$k5�;@��(,[��14����J������:�(�M�)G�#�АV�B���8���	oE���y�\����g�Sq"j|JG�	�@3RYo�:�g	fEUeO�)OW�ʃkʱ�DS��Њ�����Ӑ�GG �%WER>���^/�pK��h�LWfY�e�%���?�b����-}���A�a�����zAe�h����! 6��ݍ`s�s��Ƕ�̦�����n�Y��p^<�B��'6�:7yt�)α�GGq��}ٶf��z���fg�*��!%����X��/:̾�R���̢��f�t0��r�V�����&�I�:����z�dN�0.>&_g���O{)��c�Ip�l�ަ�B�1T��R9~���8:�'T��wf�,o��F�M�߫��'��A�֩�tl,���1��{MGnn, y^^�`����#}�׏�`��y����l�.W�khJF48l�����\\�?.�b9o����A�;�����	8n�^�����j��)�4/��R�^��Xji���U�	H�y��>����,P(S�����><��{e��}���wv��N�6���f�5�ݮ���O!�}B�)s o�R�o���n�o��i�]��JM�
����Y����U���'�`۱��gqO�u�m%��>���5�Z�� EC`x�v���ό2䴱����:��{�h�d�ٰ,?��)`��r	����A�G��em���#�\<N��#�<?Cl=~=���4� �uDy�s�}|&����1�l�W���Z���'��/槣��[�@k���5eqV��u�b���O��բh�w�����&�:����j��+đIغ"d<M�/�c�!��P���:l2DN:��,�j�L���v��|o9)��T5C��������i�y��4Ij����v����x% �Y���sf�ݵd�Ð��Ѯ����`��Sl���{N׍���PR~'�F���C����cC�W!Hh-Q�~����x����`��鬾n,��ťF��P��<ֆ,B,��E���ڗ/��8�k��{��1W@��F�X�Z{��������4��l����[�Z9��X�~M�b^�}-��<��'�;�7�:��O�<��k}��B8��m:%e�����\��Qj���o��� 5łw4��f����4�P�}��|���]��GT��{1Le%��X��X<UNx�5���!A����/����(J��y����|�"�5�2鸆�n]���$/�s54�o�Z{��ۺ�.���G�o�Y�c�X[-�\��py��ZX��c �0�mR���o�`ܦ�ϻA5I��u��9lOj��O��v$���/ݑ0�g��1���!v.��������k�h4��p������L�(�L�]Q��CE��}M��k(�=�cwX�n��:���}W\�_I�,���R����Mm��I�v�&��@8�Ҟ:�`�&27k�>H:6�XB̈́>Q�ZE�lգ-W"��|��Պ�x��&�Q������G����vޙO�鈙��ښ�%p�%�I�p�~�}��<ex�����-���ک����	;S'���s�C2��S���@�����]�։:Y���^�;�A�<��s@oݝ�����@2�g�4���\����]��]u�kL��l�v^�A"8{P��1��R�⣰�|w�_���/ޜ;e�{�f�1E�v1{U�Yp���Ô����ddLR��{[�t�3�\�Y���)�*%�����O^ݠ���X*�F6���	R���5±2�e )�LJnM��3{�+�6O"_�xj���zs��{��Q��t�7׌���^��oq:�ͼq��W�E�~���O\ތ�ǂ�����-����6���d�PV�%� z�z3�1�b�����	�kk+��~�-w^��2a�?��wE���v�"�����(G�4c�I=i2~���d4���1K�l��Xk�m˱q���ON�xh�2O0�_C�?U���bw�k\e٠�����o����'�
r]R��dx���bA�
VO��G2����N	���� ��ss3�=r�V$Q?���w���/��W�c&!���;�eFjFB_b��P\�K4�z~P��w�^����;�	,k��M�0�m�B�0���-�e����I��4"�b����xu��֮b�~T;B�o�n��F������3^��]��ݛ'�ڿ4�ԓF�≙n�oYF�lH_��r�nrp��՟N7S�Y�!..e�Y��_��Ζ��[w;>1���%�%@!I��ve�B�9P���}ߠ���Kn�L�3�=��FԸ����=o|W����[�Ҧ2���g�_�t6�@� "B�K�����y�����{��{��M��m߈�ea`7њ$TOL ��5|����}���B�:�Z�.y�a�t�>"�ʕ��
��>>Rͥ��XS�߬r0=��И�T������[)V�j_��o$z�Q���q�����oH� '<fF���d�w4�V�CŐx�qJ_;|oV?��y�\yo�λ����@���L¿��+$��tZX�����d�CZ�u�3h���*W;Q���T<@�4�o�z�M��VU�`ef�q��
��'v�X����.r��z�A}�.W*\�c��Ј��۶�(:�Y�v����h��;�_��ɆN8)0���d/
�thyt<�O^ؔ]Ԡ�so��m(htU�J�*j�T�%��K�YQ�T��E+n�/�V�Xq�]}�f�)���� H���5~�xh�4	�ǧ�h0�ģ�8�P���Jf�T
�J�Α�Gk>gpdC�����	ŕ9����G�u̾�<-OHBB�g�v�V �pӲ����5�'�歕�E����i���-,�v�*��qm�Vc)��YF��u*�Pjݷ��&�V��(�()�%���(x���iF���Wʷ�߶Q%���N�Q�۰)V�]�9j�O�%��R�Y�=~��2��)r����"����B�72l|���s^���\<�{HZ��&TZ8 ?�H����v���6��}�#w�i� &pO��,-�ߦB\��;A܊��k/l,y��'��:Y���[2��Tq�<�7�=�e1�0k�뛲vBd/bT/�ǮV}!��O�uԏN������yp�rձ�$�=�r> ��3��ȼ���Hjw��h%t�G�vt��KLo>N^�L�����8���{�a0�L�+#Kp�;b��a��sU��Φ���7tP�����Wm���Uj�� �?O¤)Mg�9,�4��F'�u��[\���0TS�/W�O���a[�0ػ(�z��|��\�Ŵ���5�(���`��r����ژ[!z�����bp,��zI�P�J1qLM���r��u�귣�Yw�Φ��1�yO��  �.x��g���A��q2�o�u��&������B���=̷������#�+�+�S�wK�t�{�e������b=ac�	323��/� �S)��нt���{��y�1I]!8.��^Tc�<E�)��|�ꊻaz�5.vP�A��cp��L����g;.�tܶw�?�mL��v�R�����:�����{�����$v����Q䢪�;-�v��Fz�%��|��Of��.�V%�V�/���0t��P��*^��h_+*'T�8ˏ�qu��.����x1_ΨW�8�߳HA|�x\��mĜ�Ɋ����fW�.GGk/�g��8�j��{I�~@"�d߱�C���.$ҹ��q{���bZN�;�/쉼x�8�r�Z��%����YS��V�����&��<v܏����Zt���ܷ[��	�DPk$n
��D��.�� z3��Y��%���J)h��֣�K�K�ŋhy�n^�������|�c����w�2՟K�g!�f��ЧD8�;��be�����I���x�����CO�2�|��^�Ѧti^��a.A6�2�:��US���^ɖ ��S�hG����龜��O�/�~����Pb1��I��8^���z³Iwß���-�l2S��.�$�$�)����6�����n��R2��'n�;�z[_y~/�<��Ėe�=��׻h��/���yf+a�O�\�U�+L�P��T�
ʻ�?FYHkwk�m��It�g[������t�!is��R����M�<��[}�3�Y�O<�;�����X��C��7��KK����c۶��fcӐ�L�Դ��~Y� �/%���Y�-�v�]q3������z��/���^��	A�4���;v��owq=q`�aht^�n�gygɀ�qٹ����'�&�����ީb�H؋K�ÚG-�
־�1${Yi�Oe���Y�^38&Ѣ���zVń���=�{�t���fS�iT�hO~�H�e���J�aQ<�*	u�}ы��O��4���	$*�3��]��M棌�'�tj}�3ro�ɊG�ݩ�I!}�b;�֌�,�?��S.�X���B^Hg �ubZ��QC�4V����
�,P��q�i��d0�nh�����}���GU<�MB�^i6��%B5/��9�Y�����^��.����}<[����q�A:&D�m5�cJ1޾�V�6B�I� �P��;fc#ҥUOL��/����2Ƣ��ǋ��:��p}��5��SS�#������q�ˑ y���Vȿ���G���nY]L���#%~F��+�C�0�n���'�j�S$��Q��C��*6�^�}�0D�3��۫WP�6�ar/���}�f�$���%����	~L@�ג�B�Ĉ���;�;�[����w��E�"�D�ѣw!"���{�=z'��[��F/c�}��������-���Y{���>�L�z�	ŭ{6��.?��R͐f3j�(�4�\�����XtP
2������q+30p�"R���,=��R����LѮ�ZY�T��ʿV.{��8Y���_������d�n=��[�f\��ֿ�l� ��צ���Ƒ�9�ƽ2�h�NW���ȹ���n��JW�,>)<oǛ?�{m��feK<+cb�nB�_�38���m1,�Y~��Gn�a�{KⰐRF�'曞������3v�'���&�JmseS?����r��ɏU��Ķp}/&d�[JԸ#[�=5�dzWfF�=>��42(���ڨUd��9�����ӻD�M�K��ۂ$C�he�N�g�L�`U�=�ȏ���끠�ga��~�EY�E�݊���`���ۯ��t[�����d\ĉtoe��K��/=�B^n�7��� O4�O�Nh`{����B������%Ո�3��J�Q��La��Jg��o�L���|M/�}�\�G5����NNƒ�� ���t�*�|U�μ�1;&�uM���Vs�l�g����N5����1`���B�z4 <8^��\$o,.�z���wk&��z�'�_�[���P�z�R{�<����u���[n��U��ˏGl�v����I}�i�y�t^g�lp�Jz,��Ĩ�����Ϟ5��=�nsv��|���x�CJ7�Z�%$�"�ȁU5��4T�g����@��[�H��p�PH( ]�!0�E#�l���eY9�b����m���WX�ԩ� n�������7�z]�#4v����~��4Tuass�ig|VE˟Dl�_���n�����]�r\��n�����t<���BC;7pGS�4���|݈�S�N�HĂ#�#68�)�ڐWSE�E���b�J��K������c ��
��������6��d��H�9�B�Ĩ-�q��.���tI��kf"2l�te�G�A���"��i�Uj����29�V0�+C���!��&���&R�gMLLp!|H��D�68<.��z�iCd����Q��Y�h?�/o�n�9��{��$��(L ���3b�\֢7\Hf���ڦvE��e8��G<�� y�ҋ�ǻ��SX�eH�d-IA��yeͬ��2,����#WS">C�v�Uho;�}H�bUC�T	�e�h�拴��Ԛ�.փJ�U�4�o�+u�=�pk��@�^�%n�)c�5�pl�n�"(�n@�%���sj�(,�tu\)���
��[i�����������3��y�j�W�b
�P��op�8�m�"�r���v0�*����T��?�p��\���|�}��P=O���c�����D���^1+f�����}�?�v���4������ٵ��}ruРi�BE�cD���rSx�db�k%zsY[i���^��6õ��4KϠ���V��sł�ym4��D��v���H�T,��E�(�V�4�Z��ش46���s�~3F�,k*��^s< ��'�&!!��keOeUdx���eW��\�rQ�]I�?=y�?��b��o	
n/��t�fT���7^{��T�T�jN�Q'�4@��q�����`rH�1�_f�����Lv*3�- 0�឵)�q�@��֓\�1��q��ZV�M�����eVsᔑÔ��՚��X�v�DĜ�y��gdv�n?�*�I��d|�vv�~9�lXx�s@L���ͤ'9$�M�5��Hз�])U��uA�6#���Mo$q��,�;��sʇ�.�ί�ƀ��O_7��`��6����@�h�6��g���[��T#��>��x�]�vx#
���߼@w�K�Wgu��7��K�vu(*�f�_�7�o��?`�b�%m��%�C�W_��-^�gs���胏t�-u���o��rB��T��sƋ�qUʋ�}����Y�����e�O�@��H,3�՘o9�����Q����+jM���=��v¸U�V�N#�O1E�qw�w����}�	��-=<���r��n+6I���^�s���W��I���&��H�lOd�?���Y�9R)*`�艸�b�*��P�=�i��l�LN���B��I�)�YM��[�]�I�-����ڦq�Ux�e�z�|�'+%p��P������4����\��oД��lLc�Ot1(��CI�X,`�x]�.�ۺ�?��+	��4�?����TE���s勵�0d�D�[r�`�����o=tv!�Jm�Z�~�~gE*婏5��j>�|
�]yj;ln�_`8Ϙ��;����n�F"�W�t��(�-i�1��l�jBU?Ł��l��3t�}_���h�*�����R�$��ɐ�-�z��+4����|H?���mD��n-���Ǣ�%����31*���6�vb;�kb�Lۈ�-�����e�������\_Z�촗�c[��I	�����&K��@���C�3�\_�i��dҜ����:[m��uI���50�6v�( y.�h�rٵ��A����ӥG w�	��I��V�_u��|��  ���h��(ea�#�C�ɱ��)C��F�Tz��Һ����ֽ@�h����
�'~�/e*{k?ҡ2�B���S/[@=��~܏~��2)�^������4c��,Z���#M&�d�ճ��A��HNw(��c��J"�}��r�����A�FC[[�j1�`�F-g;�8����?Ɂ=�_��nZ�����҅$�F����r��d(?�Y��ډn�֩gA��ԇ�䷌�;=�J��S�'���:v���0-JSo����~���������������I9�2�cC�u��G:q�}n�Is�nO�l����5�J#�Ȅ��F|8gɇs>\�*�~>��&p]klo�"����I�Gƺ]�q=�ʃ�����vC�D���s��Ƶ� $ �S�� ����B�B'�bj32P��F)�eD�ì�g-�wv���>F7�U��G �Y-zn6�<����0��[��#{�>���Z/V�A���o�B�:�Z��鿹��R՘���:�)�m�P����5�����O��5�����^��I���a�,��VJ8ո��
�b��J,(�y�������J�V�����ż��6�)F��H߄��4x��J�$��?��o�y�(=m���f`�^w�>:���b�BwD|~ ��A]P_���, y����V9SkGA/������0�Ӽ���È�Qw�+>P澠��� �8]�U��x���T�L�����i�oX�N-����������`�.��0���k[���'��O���.=�~5��������=�md���Q�U-��y�_�ʵ�h
BJ�6�=n)D�G�Yq7		�ns�}y$�I994�x��)e" ݝ����q�����ɱ�ѭA�#���gjb�uE�M���ۺ.�dBP�#�[��S�:����h�fO9;�$�w�]&No�ѹs�:�9�?�j3�I���[Ѽ�����C������&w|���X��4�w�ݳ�i{%WIwoN����[��}n	�?
�Xl��iOt�4�>�{_���f��؜��������24��a�5���|��e2����pL���!�)9ws~�M$QJ�VO<�@���q#�d�'=��X��bΚN��Y5H�����I1F~Ό�x�K��Y��-sX�8�KD[\p�G�X?�i��NH�/��uH�ʿp5*���{k����ZZ�l2"�Q��s��$��|�g&~x^�W��5���SXID��]6��7��� ��㒹�D	>�P_�|Z�0�|��^���E�8u��X�]@k@v\�l�ȗ�:����U u�2�Xw_9ġk6N
S��`��Ñ7�wwv�l�S�k�'��3³�s�k����+g{p���qk�N�ұ|���B����U���f&��蝧�~Qق��p�&�&h�p�
ם"]�����0��!f��'��d���5����Qː!�՞���9c��'OwQ<:�:o���z����ٹ�(9� h���K�ګ/~k��%c_H��+�?�\L$��%�Ӹ�`֍-mb�"#.3��f��;��ll-�Pb���~!�>�3���È3o&\�㗸V�X�-�o���eLvr��.F � ��IO������B2�7ݡ���";��|���z��
l7��򚵂6p���}���V��?)��D< b�\��:}4ҨdN?��	�*���L�K~��h�o��	61.v�4 ��� X"Q[��n}��K�:�?��^��zR�\��D����6O^B�AM5U�)�,P��)�T�Q�劜�NJ�n�Ϡ��`i��������4/���啨��]z��a��� D
�;��IQ�P�a��%h\��Iۈ�o��� �4�n=���y9x��kva�u�M�� �Q�އw����+�r��X����e�l�:�`���~�a��AV���	H6�he.@���>stw�^���o#FE��K+a����;�&�_HW�[�ܪ*�����2"�W�P&	LT2/�/kg�N����L������H�������D��T4�v,)��B��Ue<�+=�����޹��%��^HMd`d��S�0�?�ʂ6��h��y��T��ʝtk������uQ�c�v`$�-ٟ�O`�fP	)���(���Y�|)������!"�dp�F5>���]� �m�K��߄'ʰ�v�����a5P����`O5����/ҷs�S5��M�r;d�+6H�(���v�0Qx�]3v*]�Ov��SUX���+�En���c�%B���}Vh�rb��ڭ<�' �T���⁛�ҵw�AF�M=g߳7�.��y���D\�}*A�##������/��O�V����-��z�E�E)9��m1�+�1��`�v�F7������+�Mcc.�,N�rDY��
:��5Ʀ���8�x�,�7�̒�9�|���,�OǍ�EEE뼳�+�m9( ���-<��Tm�`6�~�:sN	�Q��ڵe���r�Ly��pm�c)�E>�lr?'�=�o4_��H��a�ʜ��l#�)�*d �7ӵ�Y)e�Z�v_p�i:�rH"�.kH��~���]1WX�|g��NI�	�̢w��S�Wr���oc'e)�x�[�*;B�6�,�y���DH��mIm���#�{������T�k���T�>'��Y�4�{��15PۤE��ҷ�~_�������Q�+Sg��fS�L!U-OC����1�D2(曢�L��7�����iL��u?<��i��6�R���:�hJ�Jګ�0^���AH�6�
�C�`JCkHx^t�Z��OM�b���Ѭm�C}�/ck5F[���3�t+�<��}
[�5��Wn���_��ZO0��H$��W�l]爹p������b�񢹟msmV�n,ck}�,c��ײ�<���Q"�O���ta�"�c|�/��(�D���Ϟ"z��x9�[�o�!�iu�wXX-��Ӑ�����e�k�oCεr���{������dܳ�?���B��P�sT'�:i[zQ0�տs�\��*e��9J�A֦N���GY9�S/R�>h���w��qx�j�M�dC�
�n�������qe�$|S�Y�5���_�So��	6}��{5��䰖�br�ӝZ��?� �_FD�3g׾�]4瘜�Cש,mE]DR&��8%-��j�܊�m�����sp��CW,
5�J�Z�)'�ͭ~tP�/�k��;Bޝ�����-�)+�z��T�����-Z5����#/M��K�JWf`������g�z��K���_췮K~���4�i�9ih�������# ������8���ZK��#}���}��CB�>O�v!(|�(e
�@Шe}[��)�y}ޤϠ�"�?�d�\��Ǭ�)�'�p[_z�@�X����;5|+��ʜU�W��y�M���'�e0��{�>�j�(�?v���&����֪E�R�R}���T@�t��R�B����e2.%J��A�2��,�XJ��,�Z�.�o4MR2�������R�!���G��]��M�Wj=�Jl���6�]$�7}�'H�4bԖXR�[a�X{Nh:	L���AW�4G�4x{xE/fS���Z�ڣ��ipØwPYڮ�*~���l�M��c$~�D�XO�;ZKÄ�9&���z�J��q�	_��.܉h���0���а�j��-"A�!vqܹ�q�P}��|�+�<�s#�_M�}
>�9nɉ�2�^4�Q���,g�G�����H�ո����.x~8�o?�k��4�JE�
�R�2>'���u������0?��$| ��R�_2a�BU0������.vZ/�u}Єe8@�O���O;k��G��?=�}�w��	�h3ř�w>�	h1�KC���4�7��-��q|t1�!���w��[u�����ཟ�%������2f��(�{��b'X��N�˵�-�x�b+c̸��H��,�\t�6P/>.��W�kf�>�3���|\s$��g�g:(�0v$I���@Ov��5I%TfՆ�Oz���^���xws@�'�|���e�W�B���P���X�� ��$���]s��?SUIJ�.1��%���X�,Z�\���x �y(��F�`�WVz�|W�Ÿy�7+�/9�n��j)i>��t�݄h�w�TZ~Ͻ��Ѧ�w���?�Ȍ��ޚ�i�&�-Ɯ}�'�ݠ}Y~+��z%k����_��B+�I�R�+	|ph	�9�䋌C�l�@�N^�\>�X�p8�o�z��D@�ƝT��T�������0�`!u4rβekC�6�P��w�	�L���ս͸���Ƞ%��y-�OB� ��`�ѡ�-��n��2��v�V�克��xc��ϔ��=S�?\��B���61��V�zvQ�q¹x��oL����tG�I��-^r�����F��H�e�G+N��Vw!I�YzϷ��76���S���� �(DQ<_�圁��Ӌ�bf�P[�D:Y� Qo;;���FcR>�һ�
�njA��f�fK3S���84t�>s+���$�<�������w*�n8/�~��b� _���K`�*T��=+D��$�tm�HC���x�\�;��F���~ya�B�,����-v��Y/�r��z	��{�9��׈E���q�Df�=���B�Ɛ ;Na��B0����kA;	\��?Xm�]>�� �2<�]��ą���c�LI���H��ľ^�����r!a��W�.��$k�8��AiY����x��d�.�TDeV�!�����율�o��S!;�� �_�|ꆚeJ
�+�ѱZ9l�_x�b�����S}'��<�����B�H|��u�G9�����;��X�?]�*���jy�'Z#��s��F|MzS���y,�.�j�Ԩ�r��C>'��Yb��0���ۏ�闏�/�����~�
Z�J���+|���������	!f�J��q��=[�.��#���!�����A�|�> �8��C��f2�gZU��$W���-�7U�.[S��з�k�N��t�����" lkT=����cM����~� ���AHh_���F��,��ZzN����c���ٚ�:���_�ݖC���xX/QG���������n��EE�����F�ꑿ�:�'��I��+:��.�|��=�����/��Z �h|���ى,���|�Z��7��7Ue�}��4�<��N��}�z��_���E���9d8� ݍХM2x���#&W,������Ai�?>�Q�ώ�=��&6���
�V�._��_b4v���d��k��5��S�"�޹{�d߀ف��d�
`��)Fj�i~zr4Ƹ
�1�ݷSƙ(������O�Bd�s��nB�c��"�X�O�lTE{���+i�*IV�\�����_�7�ͧ!�� ϸh�/n�X���͗G��u���Z:!2{��Ih�@���A��������D�o�vç��� �6.c��?q�'�Xtp>����Zε�(��M�X��J��V�QZ����r��&%X�)ɕĸ3f��~�/����������d�N��wך �y�+;*vb�r�2�M	�|v��Q�|����R�^p?Y-�P�6F��JY���!~\Ր6�>HÕ`��l���4uJ���Fv�'�r'5���nz�a�O�ō��R[��������W�L�3�ZV#8R�$�ָh�j�T���:�q���{Թ�y�r���K���_3���礦vLh��y��Vt��.SJ�� �4��"�DЅ��a?���2LJVS��W'V�p|�z~oA/4A�S$J)��h��.0V�Yh䊟�Wq�dO�F;��8W:�a��=/�`���\s秢,�fW�v�	�e�{��@19�ZE�Jc���Q�i<xV���띶wvQl����/�^����\Hy�@^��V�Q���j߼W��㧳�M���V�oSh��T�/#\ͼ˘Z�E����c\}�׈h�����ݻ��UN��0��Y��� ��Xl疷q�X��o��;�	��s� +RtǠő;�D�z�(�hs��b$&i���XY$����T��}��ئ6��O�Μg0M�5�}$��N.���0��ߘ!�j�)G�������������j�ڶ�LeMW�E�ܾ��鍾TP��f+��;I����E�>�Є���-�E�a�������W<��gs:t�-�%r@[4g����' ��ʙQ�qk�'k��Wj��������b�m"Z�j�b������f�p_���{.�	]5�v$ǣZuv u�)�-�*~�����ܚ韜v�'W�M�w�4_���d#Vl ���B-d�-��6A�}���n�������ߢ�)㼖�Q�k��}�^WEQ���h��c� '���Á�6�j�����~Z�+rN�Y�W�Qywv��-��w�)� �֗^7��3j�C����52 �^!5�
qG�	����������{M�3�²�7S�K�$E,U�Γ��{�0EHn������N,�W���c>�~�my�Uل��7UvZT1��у����jRy�9� � ����0��ΦCZ+X��B�\.�+/�k�E\�$/;��Sq�_A��O�h����f�tX�bmYo,�Cx�qgj��+f�</��p�ĘZȧ3����h#���Yw���gZ<�q�����)���Os*�g�)������֜���5�ף�P☰R-'�h��7�d���s#�؊z���)�u��1`���k7#w����g}��K�f�Q�'M�3c�b+MՅ�H���.�R��o��3�����0��V~�7aK0#�P!��Jd6�$cPj�ġ�P"ɩz����?���{�+�E0�z���a{�-�!�pI��Q<�%�?�m��U��+("�+�����|6��"�����:�����U�9\�6��ߦ��b=l�t�a�ә����8E��\1��#�$0vp>m/��~[{m�I�d���g,ݝ�}���p���ݭ��U~����vۯ��H)��;ۦ��[��F�+�k���:v��N��2-Rƛ�����+�j8�ό����Zdה�G���>��0�Z�'�ɝup��V��{�$�B�?�ep~rx�,cb1jюr��W!#{��=�jd��xM�,{B?~��D�tFW���g���co~���m�vmp_���Ђ�u|�o{�^	_���4 ��m���l'�2..�Z�U���W<{������y�Y�-c�oa�Y���q1�j]z�#��.��ƙνJ(�͟,!Ͼ�[��>�:SDW�h&���<�^���X����/����r�̡0>�������Dم�ڃ�=[ �<k�?$wS߾�Ly<�\�t_�>�#�}����gC�4���ю�,B-l���� ���MG���)�D��9��?�-S/X<��n��& �S|ۺ��6�����
433����N��<���vq*&eH�B������G)��!I�]Q�er�ڨ&J^�M���3�7�ewL�ٚ��t�1��w&1��-�$��{
�5ބ�ym��f��	���S.s� �yY>�xOu-��=+쇳��]�Ęï�tE=X��/i�#���U]�gJ���g��{�~�k]X{�Q��sYa�iJ��^�&�B:蚦g��k��!�F[X���K��q�<�aܪ�A�^f�g�5���G�������i�6��"U%`��'��u��蹵�+I�I�s
�����@�y�F5��-�T�t������k�rO@?���qyM�U���e���F��P8�S,�h�52��MzAc�5]����(˻@����BӅ�dh���D��6���y#r����)������(�*�>�vs�!bV��w����Bu�p����`Z��"�kf�9dx�D�Q$y$u*7��f΋����E�k+(�x�8�t�h�*��V��h�?Y���c�;����$yeV��B��j�i���Y�^�;�h�j�o�n�V�liޮ1q})��
ʇ�zm&�]����Ō{�y��+q��N�-�=Fz�)/�q����k���ȍ��>�q-#UK$}����|�fNkk?�֜匼=�O<�vU��۾RbwP�Wl<�HE�PG��ߏ�S~Q�#cףtLf�1���F-�\�7��K
�sU*�F�{j=Ł�ؔ��.1������G��$?&����'�b�o'�Z���z��6�����[Ѩ��~�n�@4�ܱf&��Ѧ`��?�0��wNEoyq�әU���v�[<\O!��q�7�U�(���p��_�#9t\�#�VR��r0��⨻����З�)������s���S��������uQo�������Ep�6�wm�2�v1�R� Tf<�q�k����9l񳫆�RJx6E8��s�ra���b�\H9L�y�cQT�u~��N�݉������*�9p�
l�I!�K�-S��q�hق��et�4l�Ҏ�����>��4�Mcщ�~�����R�G�ti��ݼ����u�V���_ż���A3�oe���Y%�5�5���i;�\�j�7E�G�";�����Rߝ�����v���\��֓?np��;��dv��k��B/߂�&_Yu��y.Gql;���߶�Qʳ�/�g�OEhS\���F�N��\M�1�e~;���2�g�k��#JJ_G-Cjʱ�4�/��~.�;J"�g1�hz��$c��J}L�:�o�a�b��NTYy�qL5*_#��� �c���Q9Yq'y�ǢhV�,�ϰ��S�� ��g�oy�(#3��w�9���v���E�s����=ǉ_h��N4E��D������yF>�����.��$Ei�Ntv��E �K���{4~� 0�T2�k��x�C��[�ĩM�0N�ߡn�3���3�;��e ���� >å�#�_}��dr�ᮖ��He�FEDR�)]�����޺�)��-�	B�+[��hֲ�̿ �Z��T,�����e�b�.�0�-)ꥃ�fk�ʜ6t8�9���*33��������`�H/YmW�Q�y_���n!�KϚ�~SJێPR}!k�O��MU��s�+r4��待��5���:��i���͡���t��^��W���\|y�u<�'4-��Xu��gF�ݲ�?����?XZ�C�`	�kC@.�w�4��s�%%��������8J���߬�žMp��hԶ/���ۆPh�;��V�I	pb��Y"l��k����|ƨ�<�pe���5��cDX~^�����!'��3����l��:@"���rؑ�|
�D˟jg��5��oXI�ڏ�38=}�W���%6�%�n��d޴7΅���ϞL�j��������,�mV��,N�lj�a�g�g�b@���3�M��Lj�K��Tm�>�\PO�0Y<I��[g�b5�pC��l����W��γ�Y�EQ�����o���/���9�2������������	
�Ʀ�
d����M�������:����5����$��� �/�>R�T�ʬ΃s������`K՞����a�0����}_�N�i��#��q��J��j&���`!����?`nF��l��
��N�4n)A*�@�,#X$7r����y-��;ڼm��Ͽ�Qn�|�4C�D��q��>C�R������Y1%���{=��NQ��=�&�G��Hs/e�oCD�"���t��dY�@�����o���q�L��!ô�&)�d��$��Z��O>J;���j�%?�V�2���WK�G}��39U�$b���7��J�K;��3�*J���0���d���0����ѧ���ҔUɣ�|3��Qӧk�=�J1�a����b��kM�>Nۣt�35@�*��a%4���R�?�j��o�b��қL#ۓ��"��\��Xr����
���=n>O��?Ua�[~z��������A���?&�����"v�5.Q���iGgaL��9B�֣��������������ڙ� 9��ICߢǜ�A��u�;�{9�[A�����%��_S��l�Q`�~��<��~@ŐP^������ރ�|�>�-���0]j�V":J�>�1�D=�����zcWi��J*ɢ�?ev8��x�Ȟ� �܋��~7��CţTv]w��ǼBufrR�3݊$�:�{ު���%\V�Hx��>�O��`�W� �Fy��3�t�+v�r���^1�V�X�=�������K3��ip����9BNhJWo��<�
��̇)����;�\��~�I��ʇ����)�,�S�F<oob���T?{~�B.#�r���U�d�͎	G��y.궸F��IR��C���e}�nt�T�y�b^�̪�I���x�H!�u����+�U�t��h>I��5Z������U3}kQ�"�r�*@VL������4x�-��v�ٳkK�*Z��F'5��g�~ɟ�UZ}�B�%��lKx��^ϒ'T�k����%nDK-��:��X�4NK�#5{%2���J����D��-3/�{N
�g茒�s(��Z^qMv�;����Wq�7f���r�V�27��ˤ�_�뙮����<��Ԫ���<BR�H>�w��VP�����L���{�.���e���f�'������a;-��+�}���|s�
�AVwg,�4�
���b���bn�*�m�)�~AՅ�2)�\��1�61�޺���z0CE)'����X<��>���`/��i=.ģ��tSn����8w�t���Dx�'���%��*�շ�n�i����2��8�Ü���V��D�
��n]1��V"6��i�om�!/�[��.�JI�)yn��v�2��iQX�?��mV��L��G��J���p3iS�c����xw2H姄D6��Y��]#��KVB�Ҡ^LSxrày�uD��.�L�������ݫ�ے��MLx�!�k%��%Էy�)�ft��bFxChVƪHG�K��dr����8�Q�a�K�J+��2 ��_sq���;d��gޙ���r<W����eO���pEI��>�b�آp�ĉ�mW���(K^���Yݴbҵ+1~pL�c^�{ʫZ>c�'��?n������v�=��4�DHJ�֐�a��Ji+��nZK�_�g��������BAm��_����~7�F���)m�>M��+0GNӨ$�����VN�.4/������oWV������kCj=#����E�.�!T-N�{�Z��E�Z':��������.���ǅ���%gh�%H����,*��D��8�}�����K���� ��S|�o@�B�ʔ�c���i&0e
й;�1~��;.�&�*��^��}s$�;	�P3wr)+�0]�g��IZ4�s�Tkxz���ϭN��������c�[����p�8w߷�
Y���]h���4����I�J���hգNك��i�I�������G"�6��2�ߵ��=��7��e�����W�B��0�9��7;�x!J���QH3a�K�	�NR���G�P������o/��D��$�)��=�L/,Z1ʕ��(Kۈ��(C�7����HD�=«P��85���9���VU)�j̮��&1� ��j����FCo[~
n0>s��������v�dq�ܻu�Q�N�AP��7��
������ybب!��[�8�&*h�d7�5�ػ5�!�gL��z)�ϸfx�#�]��5lԪ>���W�[y��M^�-/�������\\��y������-V�v����>D����,'^Y�omܦ��UzVa�~$R�Plf�DA�$p��#��k@��}3!|���#�>n@���S�Z$'ٷV��(z���TJ��@����]�	r�w�gM�*#�`2���~���B)�Ce��5V��nZҢouY/��t
�gn��>���Q����������G�Pأ)���vz:\�M-�Vs�u�;����N�j��a�ۈڅ����A�V_�M����V�cة�hZ �o9��݂�H��RXg��$(�41���rz�Q��C� ��~��G�KK7�2_��9��sLN��7)�y�H��c��7��wC������yao�خ���$k��y(Ę�Zߏ�M��g ³�#7�=c���o	��5#�͎��a���5�6L7�hk�k��WX~�����Y�3qgm2>�0�ؙ���!y����u�83֌68��o��{���6,D�L��r$��|�< U�|���
Q�!�>�7�G:����į�>;��,y֤ăX��r���j��4��ΰ�����TV0�~#��^�+���k=]�hoԋG���f@&���J���eԔ�h�=����~5��O.��ᐼe��1^��y#m�H�{���N��Ѐ	�P�����	�U���B����\�3L��Z)>,���眏W��%�Q^+��X��������k�V���̄����$NX�q-��_�g�S�&-=*1è����%Q�ä��z{x�x1r��Q�w�l�����芡ꮌZ�y04ؗ���;��^9{�k������[����&�H`[T"9]n���\�K�o�,Q;�t��M�iY��¨�n/&��������"E�z�����;c몿 ��.H.N0��C;lM6;���Eo"�e�����|ޓ�l����o9��
�����, ;R�H�vl�[����2��;�9��g�Տ�������3�X��CCN��Q��)����5W�f�>��ǩ�	�Fi�$YG_��C��s��BQ�,�v>�w��)g�_s*U ���aΝ��:�/�S/��^^�NY�;4���g�,;���
�m.NR�K[O#�� ���>KO�Y�];�Ӟ0�l&ȹ�g
���Y:P��<��^E<�H9i5���4����������~�E���[wQ2��7љg���n�υ��͸L`M��7�-��?���&8+���o/�0�d3r��3��̓K�_���'�y�ˠ���x��v���rl��s��O����ވb%�!�B���w�CPB˲��/U�q���܈.�dTS��RWbՠ��._�u��9w�͵d=�J�i>��p=��4��4�<Oȹ5�G���$`�<�$zjl�gQ�����q{9���ʉ��M�3���!VG�t%�Jԋ�K�%�7"�o�ká�'��֯�*Q�~`��[���[�p�H
bU�_?���\+Iu�Y!����4}굶�<� r����z�8吤爋U ��3���ڍ9O�#�6�>F���A� �=1�`�^�cxV�0�ү�մ�QD��ȑ��P� ɢ��.��o��vL��0ߓC7�J?5�BC:��x��>$��c�|��>��Cβ���?c�U5!p�N���B��ܜ�[$�W�W��?��ۢy��I��;r��̆8��k�7�uD������}1Z���"��9�1�O��sMa�� ��zz�&\4=%�A�H��1O����������^�z��߄[�k�2ȿT�C$G�N����֋�J1W%�qՇ���*�FvP�Q#'�r��
~Y~,R�#��;�C֍Σ�sR���H%����=��`)h�Qf�,N?�Z��_'{�/2�냝��̂o��f�O����q��Ak��"}���/6���X���R�}�"�of�Gz�����S6�I@#�\��K˽~�I헕6b�=�/G��JpTX��וk_WnI<�,�+�o��$�sYQK=����,�F%���u�x\��s���� ;kB����ny�em���^\ y�!�Z���U+c��z=��P����~��Kh$����֒Әf��%L��?Ը8�i�6�o���w#�	c|8�Xw)�'��7yE���H���&��w�%)��,�N���2��!\w��P�]Kv�����%���͍%NK��l#vQV�Q-�N��0����p�\�T~���z뇦��{X�iF���[�n�Na�]#JH��tw��1P����F7_�����/�p�s�s���3�"�� N�{.���nP��G D|��I��4MX��k��~�F�vo�<ϧ$y_���Ud�ԦX��V�М���4���5�>eE��Q�u=�H�f�Ņy��k@��f���I��T)Ѱ��{��X���ё�M|u�Y���M��	ay�è�/�˙#���=[���X�.�h�K���j�U"V_��.?��;jE|�X�,�0c�!�Ph̑��t�Z����#�B����<��Ӓ��>x!@�ae ��ý��%6�È����t�\��4'�7c��d�}���_����q�+A�jUU-�Vs��8G��T&���7�(j������h�|������χɹ��Zvx��ɺ�O�t��Z���� \tZ؂7�D��ᲁ/�-�����p��I겳�lJ�u{(�n}?�z��K��=��'�DbUٌ�XE
��&���p;I���P	�;$���>�R���޻��V��Ǹ��Ʀ.9
i+֌�����l&
��C���-a�u�xD�Ԣp��J9�u8�J�p���˴��W���ᷧ-Nˑ��ǣ[V=e������&`� �IkT9�yBC��*s'*j�ĝ�^�-,��*�P�I]qss�:�gu^��s���G����G���.�(ށʴ�����;�*tm�p�#o��w��P�N�ԋ�bG�)� S.e���MI;���CT�oqor���uj�15&�ɚ�]'��a𴆜&�`����`J���#4���v����������a�j���Id$W���(��"	/��½hg��>���������=zdS2��̨D��O��BBy�_|��FZ�&O�T-�x�E���=�����Df��L�&e6qStf}]��"�2�ʎ[��%�j�v\#�[�/.4�G	���TGG	{���V���FP���ӭ��1>+h�)d�e�۽���S��pt�=�`�k��&����*y��7��E��r�}����ӥX̦⅟����F���˦Di���&){ևlO�hO�QY��v��i�HP��ti}GA���	�HnM�T%� 1�9oE��0U��u%WjjZS���O���c��]M�ȳx�ߌ�����ᴌh�	c���#�v�}��/�?R��.�(I7��RQ�����2�5��*a�t�P�lL���ш�lQ��i~.�Y�c�N�l�j�U*k�ekwD����.�sc���O�:���" �[�g+�XU��沞}[���B+�י��F�p�����g���Q�;�D.��&��~i�1�����~�%����i�z�"�C(�]�[/�[>q�������	�my���)�G�<C+�:QݞYgI���y�}r� �z��3齥J���0�x��=2�u��x�wH5�8��F�><P2���w�����Q���a���!�?6�.i���b�5Ϊ�+��#�nM����`T�4�e-ί�����E^_����II8%C�E/�no�
Wj|�E#y{9{�J;�C����]��/��ݹ�21>@��tV�����8{W�/\�:÷e_��c��
? \yz��)"Q���ۣZ^I�1�7A�TO�=:��\�2��E�^���O����6�Z#',?�=4�L<�C��w?h�m�/���+���?3�f�Z�D����?/y��`;(Ҷ��w�\p��Ti �w9=M˶J��Ѽ
hȴ��U��S��L�)�'ҁ5MQ۸ah�^���Aoې��I���\dY����o�s� �W�5�!3��#�U�E�5���π��cEɜy��1_�'�m�ތ���P�����YU(`%��/�$vn�d�>���{�����[B���m��Up���������]�LϽ��/�Z�����:������B9g
�������aa9�l�U�a�+����v�)�ܲf�{�*�@����Kbާ��Y�S�4���V�EY�[�
��$^�'������36GP����n/q�7+����<J�R3�?Jҭ����v��/�}z�a�k��GV���1��|��n����Rv�^���D���a��7��lRҰ�6��z�z7�a&��q!��,��qd�N��k�2�j�//��d���*��$�������j���9���cY�z�5 �M0�f�cRE�����s�2~���t�Ƃ�X�`- Q���?��w�z�.;?��v~��v0�*6�!Z,/{&c���E,�&�c�*���F
wClT̿�²�x�n(*�,�a���F�(XC��l�nK~}�+P+�筨S�Kb^k����	h�#@�W���Ϗ��Qŵ���Y�r���SN6&�/I�S��J����h��/qT^���_��BH�����̋?�	�;k)����'zߧn��jN�x7��6�����3�]�M�v��V�X��Xݤj�l}nt�"�PN}�u4k��ELj��Cg�	�����j�#���/>(K�v��ɥOX�;<����u�j���N�cƦݪc+Y#��Y>5ya��>.隣;!���#�j̦E��H�/���v��&S
i/�����CG��<�K��L^� l�l䣞�lb&�͍狳^�~ֳ��/�̬�
\�Ȟs.:]O��G�Vn�(��ݤg��P���;��N���pj9�-ь2>�h���[׷���07=n8��@ƭ'�)Q�]D��������XOM�S�X>�q�L�M�:ڞ
��JS%����Ex����^���!���{.,���ф:ٟm��X�ퟍ�Vͺ$��-ϥ ��<s���mD�T���T r:d�_�U�Ԫ�T���+7C9d<>U
bCĞ����(���\�R��h*|z"g_��d����O���,��^O_�g�d�<1�bE�S7xL4q�U�;�׵_n�M�-^�m�lUH.L[�Oư�����O^�'P�'(���Q5��%��ίA���'ޕU���yb�s��3�Y��F~,�֓V�ew�P���n�ef��s#�>�m��m�~��tƫ��L�--6�K>nj߯��Q�܁�p�h�z{��O	B·�,q����#�?��73�+&s�n咓�]���i#F�܁dR6��t�\{��Hb>���viw���a��J�^�i��A���?-����;�/�Q(�0xs.���Z�ME��j�Ir�s ��d�Qv����~d"O�CYce/9�f(�GH���d�S�C���V�>>8^��[��n�'�b�ύl�Nz��)�n��=4�K�h�	l�~k�
�-��&�/j`�B1V��`�hn�IH��Ȯ�TvPw �
y�T�M������'Y���jw������ɷ��O�<�����]�-��r�v�9����rJB4'a�`M�����p����k�Y/�M��S�|�[=<��Fp�8�ɪ���	5�A��f��

ݢ�N�[�S�,�/V��~&�a��H$Q4�P)�7�H��4[wǬƤR�Rߵ�w�ິ�s�����xi};��VN^���K��.�eJ����~�`hl�����>�烵6��ù{����i�~�4&eX��Nl�ǂ����m��'���Z��磢a]T�ĝ�����Lə ���6��!�`h}�r����7�?JުG�Co�<���������/����J��p2�#�t}m��_0"?�-M!�;_hz~gˣ'z�Lj������E6����&�,��F9 =�*��O_��c��l~�K�N�A�J�6�1�-�V���78T�%/�ڍ4+A~��Ga�t��s�O���aFYY�z��憘ם��E:`�k�K��>:�[Ll�
#l������������i�C��{�sk����c����)��TF���0\������C�^�#�loRɛ� �xy3Yg�����ES�uÒ���^���-գ�WG��{�^���τ-`��%������f��L�Q����
���8�yK���2Lm�e��`�朾'Q�1�ֺ)�ɇ��{����95B)5�͕����;����iw�Q��Y����� `�B8��[?���Ft'�w��s��K{����[\ҕ}��D>��!�"�����S�i�}Sx�M����e�3��9�
�Ҿ��<�=�Q�;0�<Vߡ� ܚ���sa�6���m=H����n%ڄ?��a7��BS�(�
� �7MS�b��;Ӻ�i��d6��>7��̪&	9��O)}���8�zE+%},P-��\:�W,�P"Z �:�#�'M���t.�Gf�)�9�Sy� )ׇMK4c�6�����q﷟1�Y?.��lP�|"�m�\P��d��y����m�Szf{P�U���L�4����C~KF��3�(և���zH�u#0�\�{�7�v���3������2UW�)�A	��?��)V�\^������T -����f~�'���Z?5���l�|:�x�9��r��}$8f[�����G G|g��xW�BfJͯa'�޲Pd�m,+�אꖳ���u� �瘬k�W�� ���{�YF���[���!g��6�ȋҀ��]o��ω��|��:�wx������v���d�~.�O#2Yt����;�	����TU�}���r9��&�1�h�z*��M�y�n��(6k�Ղ�L��"er�iM�?8����{�S�lT��r����g?n�(���*�i�䗅%T}���e=���~.eS#[?RB�w�!�L��*G��Ӏ�S7}��d���"���e̽ ��s�)X��u΄�u��r+3�Eji-~ދr�Z ��^Bb�A�}^����B��)2�D����Y�^S**�ܒ�X���4������yT������8�Ph���+j���X;���_���L>��oc�qW������Kr�+�c_J��"5[o�j�db��7b�q��ug�6m��x�n@p

�Rv�a��ס;&�<�:n������~�xN�I	?)$�I�8޸�N�:)�'����E�úz�|m�uI�),G�ܗ�J�i�=��`�,��V��6z-;Iv��ANj�Fh�(���J��@�y(B�?f�h���p	�H��&�
P,�N>�_�ݏ��h�k��u�-=����9�7�Ϝ��5�^�x��Z��Pˇ?v/!��9�C'�s���o�d���"���y*��v&� ���i�^/V}����^��\P�k<��j�"~tC}�7&�v0�RQ2���J��t�Ni�x��K�7��[	�����ד=��8C���:�}���vKҪ� ӯG'x�Gk���# ��o��1�̸��TE.�>�:NYo�3>WN��'@�����G4���d��:��}.�>d����
������� "����1��2
���k*g�li��_C�:�� ��`��5"��c�<�%�A'���k���DI��jҥ�؇D���%�c�v��t.�c��-J�N)�e�i"�*6G\�T)�y���Yj��ѡ�HQ5�{�CϝIm-�l�sQvι��`k�Pk�P�]�b�ޡ}c���������(����)-d�$xj�����u�W��8/��&���/�ҜC��g�:�F�n�~�뎣�Ѷ������H2I����!�6��� ���`C#*0~*gq>��0ʨ�?�hg�m<N�x[��<~�eOOE�k�����?sOfϷ�K�H���E�SJbe^��m����d/�`U!���6�{ gZM���~�0��Ȉ�js����=�����'r\�i$�M����Mst+��b��"�!�WR���5l�ٻ`���3]E���PR�#�����:nD֩�O�MQ�HL]�1E���,Lk:�m{��N{Zm;�7#[7�����S*��>RDǦaeZ�}��vRrl��Sb�'7�Ah �Б�u ��%��4�ca��kD�i����6̖��g������*�`.���v6�i��غ���!5���W�<L��̏�{���s7N�&ӯ���wA5�d�`QTW��.���
����4���M�o-)��3&N~bm�{�&:��x%�'q�Bwq���);ƫh����_(M�a������Y�ȧ�3��_�?�����ԵFI��{�W���#�2]ƹ�����e֎��i���*&�-�ءFʸ�(�a꣄b�͠�_���"��[^ i��}uwƴ�鬻�'����eRo�|�O�o7tq�6�$����Ø"�j�cL�T�Ŏ�T�_��;mؙ�WA�����-!� �����N�����ǛO��5ǜ7ַ�+?����#����W��g��D�^<����uzV1�
��؍E�F>��:�&bRĖ��A���^ܟ����}/�n�@R����[��X���U�IQv�jX�I!��~���Z-��Laۚ9֗|O�෼?�E+�NM�>xpA�3�:������{ϨV��c��;�	n���-��9 V�.���wD�Vn\�.�P[I`~����ڼ\��L�j-LE�P��`z��c=;����W���X�������&���q��v��ֈ�5�jS�(c�`+�)�{�䒺�����c�����[����┝��-�͢wr ���Jȩ�4��	��. �COj�Q��P�dL��UuP��DW!R"^��8\�lŨo�Mϥ9�$����_ITCg2)�����9�ʴ��K�S�Lj�"�Oo�9�0�o�G�8�tw���B�9���y�^!?c-��b�s���"	;��l8YыF��ĢLn �a)��O�:�s!�t��!|�p��mr|�Rx&n��2��R��(	�z�<&H0~m��b$�$u��x��j�����'%�B��'{>n�������R5t^o���I	؁���{�QK��n�ϬVz{�9V*	iL����c��G!����e���t��᧍D�1/�����P3�k��k��ws���O#�4�<^���(�A��.�a�\��g���:�m��"�
9�Yh-]�=��0���pԦ�烨�6[���5���x :6s����k��o]�F��H n�6y����z&���-[`0qe��+y�S�3sO6R���������)R��H�<��-��yk��sGp��٠�֋쵘ssy�O�ή���d��^DƢ'u���ig���-�շ���Nj��уtn|o�e׿~F�j*t}1Wi/��؈a㛴��t��!�a3��>ݗ��@Xu5�*|���m/Fps���!��ٗ����E�Vf"ݯ��dgI1�6����+<Z6��Ao�̵��6oN��r��IFw���e&����t�T����W�KN���^�Ī�lX�RFDY�'�u`�lq��ܐg�*�Ų��������o��0���}M���'��l��ct%<�����a�e�uȘc]Ĺ�m�R�*u^��7�j&_�ꕎ.��5RU7+��`�<�ײ�D8��L2~P|���tw�,w����r�5Qҙ�8�pq��½|d��{[}��z���zAR�5�xTWr�R�ۉ�6��+.�f����{(���,�,6>:V����v��ԝ}k�Af���v�U�t���9'iΒ�>��ue�tN\xJ
e��`���6�ng&��s��w�CJ<Y��rZ���3�\�YZIx��A1ˉ�n�qO��R�m�_k�p��)�&�{p�������Ւ�.�|�����q9��V�ttlVx��Ma�����R;;���R�����l�;4�㎣�	�'�b�t��NSn�=�@��`i�^�7�0No�
mD�%֍ ~�x�L&�g�}�I=��{��(�� ��L�CXPL!���iw �;5W�b'������B?���N������Q�j	𖱵T��I�6��{œk�Np��/ׯ:1i�40�Ϥx�%$�x,�E��g��&��1Yy�'�Ӫ�O�g��7B^7B�Ŧ]���7=�D�:�5��w�f=<E�Pĕ�k��Dٷ��$�5E��\y����[e�65ktW@ŀ��#B�w"Ap�O�����n{~wی܅ŗh��[���D�{�Zwb���Ix_y�cpWJ2�G�"���Y��|#$�'o����;�L�\�!�<��Iൖ����w����Xs�-i���2����庫����Fƴ!���˚+�.O2�ڼ3�o�����E��P�]k$T����*����n�
�G<z�ώ��ٝ!�cWR��즧hfZ���&���6���[�Z�
�*����.��%o���ihK�b�����'?�����v(��ڳ|�uf�Gq�F]�ϝ@7�{m�����vL����<(���H�i��gJ�0f1�3�l62�X)=t�Ƙ�e��g-햡���B!�v�@?'���-�������H�>���w���V�[�[��Ŭ�J6^b.t��M�X�B;��Vuڜ�,��<;��1�c�+˯�b�%j��kC~�Tx��0D޹;�|�:%����d�\�0uP^L�MV�.�8=���l������5�.:[^y㠻J'=�aջ�y����rRŌ��SI�ւP�������fzA"3e_�'k̈5Om��]�j�h/�V��)P\Ȅe�:�/������ᙔ��hG`�1ﭸcۑAu~R|��90Nt��p1w��y�n�5�R]�mZj�z�����P�1��F�\�Gab��/���Z.��Yf��� I��
�{X���n޴(�I��[|A��>v�9��1v��
ˢ�mA����첤�M��)�2�2nχ7\7��]�����P%�fI�-���t>��м����@�CE�"~t�r�0��,Y{��v�d�yN^�6��f��V5mG�z�&�Q�'E�����v�Ā�]ҋ�%�����m_��rj|<�7W:d��>;F�}���9����1-*�[L�O�*"��a�����s�Us����JVz�Y�d���H��&��m��Ơ����k �m X���:������:K�In+�߬�>9���I@�{p�3s>_�_i��"4:RoW�VfV�L��h�4���7�)X%}��W�c�����-��3��i�kG��]E秧?DFL�����g��獐� �U����X�L�.�jp'/�
)s��;� 8|�Ѹ8
�J���2槹%bcnL�
p���U5V6�kra�}�W����/d���i����]�����%a[B���W՟��ߓZN#�4-4�!�Y�~����G�c�f�,x� ?
��F`��[�gqb���K�O�vD)��-��yS��f�^U:��ڽ��4���K+��݁om18��XӒ�"�:��.fЌ\bׄ\⇸�W��n�	h5�3Z֞�������b2�Qg��E����"b@)9Q{���f�C7���ּ��KiI&�3
�����Iu��u͊�%���<�M|t�Ա��� ��H.`|,�����b������e�˻�2��olB�����+b7�<���YĖ�[�	j��z6֜C����U=E5`���|�mmTjN��.���4W�0$������j�ܔ�Y;b\!�z��H*@1�p�*J��l�ʌY�^�m�J���J�u&��������߉$Z�rz�Q�B}�����)��i���Vn���te<�h���+��~���
���t^O�#���7��kH�����~̍�_'��3;�ڄ�?N��ʹ8��CeJ�^Ϲ߬=j��i&׵0��
3�+�+@`�63�����NyHw�k���nmk&-��D"t�ђ�� �@����0!C:�^��~��J�KP���w��1�k}�[.��10��PX#ǉ�=z&����Q�L���'o�T��a0����:�i��\Vʆϸ��0s�Z<�u�S���|6���_���I�pWk�$+`�ͯ1�#1?]~��BA@�F9O	�q s����࿬8?����Ӱ.��T�:$��NL3�w��e������� �Ǚߺ������1��l�ؑz�ws��N3�<Mhw~��{Q��LSI���B���j�d$xd�_�̉{�>�$�5�3-���uK2/zQޠ�z��(��ϏC��B�	�� ��*KhT�Z���mf&��}�����x%		c�C�F� N�O��*��#{Gќ��uTecpfb��_v|��fpK�����.u�Ht���M�ī>�q��a���6	��jA��~�-?���A�,�]Yt73����K-Jz`��{�c�rJԚ!�m;K3wD�<*�z�&ޔ��[g��&�Imc�yٝ��qw�ʟ�����J ��Φ��p�U݌^���U�v�Z[o�g�I
�����k�����X�1�v�/~�K��n���l�t���`��Y
ث �p BN���%�P���ߵ?�U+ ��������ȅ�߶_�X������$��\
Z��~0��A�Z�s�"�0^jߓ��L���])�GV�P�;b�\�c�~�^^P���u����q��Z�D����3&���=v`}.�i��B�&�U\P�3V�~�i�QU�*r����hV}c~#��Zw��k%i��k�.�#�t�[�^2�p6n�S|zr%��;����rA�f�`�+`�Lz. (.�Hfr��~�6Iy����jAVǒ�Li�CN��.ߛr@w�
�Uϴ���9>@�-����׆nVO� +;���LwP�0d{���ܡ;}�]�zb-�$�^ۡƊ�����-�?J=�YB8�BЁltF�Et�G��j�v��^�I��%lĉR�-6��K��󛑸q�z!��!ֈ��t�	X@>E�i8��kGg�Ɵ_G�Z�].`�q�M�1���F��>�~�jކ�6��=ܟ�f'�޶�WN�&��2�� Rޒv&��u�L]NB���e]p�J7�_J�`��]o�.vB5^�W=,�w'�z�Ten�Z�Cȧm=[��o뙟�}q6�n���E�Xԛ����Wcz���5�÷|3�qj��G�R�K��k�^�	�|�.Nk�K'	�Q=v�t�42�X�*~մ��gz?ߞ�q����TH\E�R6�DH�h[�ϧ.o����(�&�|���b��ǡ�t��P#�{�1�5ް�\���K�� z>�+����K�h���] S#v�Q4�I��bv��"��Ɇ�O�ë�_H�::� �q+$�!�Mh�WW�c��mh�TD�J��|PG���u�~N��w��Z����ڜ��S��"�y<�'��y=SSdrUʅs�1�4��5����8;����-u��HSAt�eU��՝��j���Zk�>\\�X�Qؤх�����Av��-@�!糳�Y���+N���S$1�e\W�W�%��"/�^�����+Q��Ҙ.P�Z��#�e�iUv�B���I�V�
�#�(鸃���.r����{�Ws�ɗ"��ݡ3� ���43��t!��֦S�z㮵���/`�9�&>���C�;��@o/�!��n�[�6)Wm*+�,̷488a�[e����O������|�XD��mw�s�VI�ʜ�e�����m��#�U�֒0��1@����`)�vW��s�i{�n'� �s�Z�����oR�W2k���J�,̐9��x��^�N7�͆�o�@���oug���m�����I�}kռt������>�֬��[��A�R���K����0��{ȏ�w��UK9D�&�+Ҏ.�*o��c��u˶�zT������0Plz�"l�C\�|��Zb��U�z�p�qIR���ŵ��i i����@՜���n��8~���닰��N�y1wW�r��P��9��Z#�U#y�L�Y���޻������V)�����G�L>q℗K�_���Q��gHF��,��Џ�ԭ�=ϦE�����`�����������_�
����:|��r�sw+/�\�l�+��9��7�3okp
|+L_�t'�����]�Q�����ɾ5TK*L�
�]U V�:F�^7�CV��a���$V�6��s�g`��q.ě+0
ś��*R�\������z�Qj^���;'��+v)�8򵐼�s(��E��������'���ʕ~Wa�����]#7s�t�me�4D@�����WY�6��2������>��CB�S�/�e����B��ۑ��;&����n��x�ݏg�/]I�	�#;�ӡ�JO@6�Xi\0��:@�N�7�Cyzc�1��n4�8友�J��O	��-Ox[C0��=!��cj����e|s}v-��M�`I)W&R���p���gחr��g���v��y4}o��T�GP���HQX8�FK��^�~��Obk�J>#�aM�y!���Z�A�,!�N�F>�Dg�;�8��e���=]��J�-���ϊ��<#�Ꮎ��r~:�������2n�e"��x}%2ʶ(%�-�?����V�����9�׳�s��\3.�po�u7��s�v�Y���8��fN	�n:�=s����4��l��F�!p|�J/���7f�y���h5Т���p(���{j<ͫ����PNRvt���@
7W~Q����2���$b���J����k 퍕���вd���_Y��V����x�X�Ulڍ(e�w͗?�3�&(�3�%9��?�}�|�E�2S��K�X�nX�C�`� 	~�'}d�N7օxz�~�n���b鄹]�S��*��e���'=�����u�-��.o6�fx՗F( �Fz��(FC�'��Oq3?�����} �Ӡ�6��"�+�/���ç��ѧ.YLLR�^hxD��D}��Ԙ��@9x_?���7�p|�ȋ����fUJ%.X���]N@O�F�.-y�E��Z�2��ʞ�-��N���Z��xh�����(vx-�7�9V�FM�>�!O�|�^�� :;o�S��-��A�O�L�~/Y﴿_�XO��YL;�^G�� ������LuJ T`K�3	P��C���OSL(˫��Mq� �0���>��4�2f����Y�)@�}-��g�+�X�(6q�u���8�*�z�
�"��n�0χM��*`��6�z1���>����ƿ��q���)s��U�2�f1���pO�d$�����<�3�2%���A쌑GX� �_X���4wk��@_�홐?H%�hfu�!�v��p�l6T���[ �z�_��}'�R/���@�[�ݹ�{�����?B�� 5�.����Kے��`��㋣׏!����24�wr#�~J^t5��R��_+}[l��]u�,����c�L�G|�޽$kB�vg�|>�K�2�G�Ӝ�+b9^U��nk:��T���C+��.����Y�O?OZt���2��v[������ ݷ^߸K��['�)ֺ�*&�����)6M�Y=#� /2��Z#}M��GU�.��F�>Y�l��-]�y"�1�y������.3�Ȱ�^@�<�>���P�r��(���V�j60���a�{:Lu�'h�~r~/�$]3���M�m+0��ڂb�M�*]�����e��bQq�8o�� �z��q�޼jy1+�Y��/��S1�N����+,T(�Nki����~��n��uIx~�q�����>�**��f�ވ�d~S7��ï�#���n���%]�۔3mAya��#�33��,��P�%,WId��E)���	���S�a�6k��=�E+~���Іgyٶئ3x�ئ��'���n�1��d��"p����v.0���x���`�����(����FYF`s)^i�P���F�(I{!%`b�W��7`�"e���L#�>�S9DI���e�,��o����p�.�*|�+a�9q��:itSd>Aϥ�Γ�2�Y|��M��<����ݥ�\*ڧ�cl_��?	�����Y.�������^o?6�M�W�"A��>��v�+�W\>#vV���=aY����^�xy&:�:s��F�wDE�Kӡ1���wl���U�9j��GaG���_H����2�p�F�q��ۅ���|N�1;+��o*��#]6��A��B���^3������M1�<��%{���f�^��������ٛG��M����(���6�=;��'�;t��9H�c�o���K�w��\���.K����d��j��jU3����v �"�4AF��;:�;�\�s�1��� ��O4�T4�`��F�V�\�և�ZUz2��o��l�	��0u���ei��I���b�;�Wgk��n�3%ϷW����ߌ9܂%�ދ�d�+���no��r� ���K����^O��=�ɲ&�؜ry�`�o���I��w_)��u6���}z{7�Q�s�1�����������n�ă|���0��D�+d]Z���A��er�Cg�����lֺ�Eb��˙�ms
�.�:���g.z�<պhG�����eG7hxv������I�+݇���O��Aj���$\��'O�3��"|��S�3_�vk��۝7m���Q�r x�o@����k���ޞ�x��s�����,�2��NzF�~�t�~t��j���M,�}���X�ӜX;�|t������~�(�^�`lA�
+�����"^�\��5"���F���E:j��X�s]]�띥���؉暑��7"F���!7~��L�;�m�K�1�)�K�\�T��*Y{��\��G�(>�Th*�#={���`t�j�=s�ڋ�%��4�d)�h���u9�o�Y<�3<F �1u)���1����>�;֕66 �	�V;�H#9�ڸq�v��Z[զC��JL�%�Ua{lI��w�20~��NOO;��̖���.}T�T`�>s�Ve�+��ɳ�.4IǗ��ߘ��mй�M�Ð�"j2"�[�jHȁ���9,υT���iE�7v�X�}EC�V,����B�.=��������#p�0�)��4��k;�vi�C@����|���o��}}o�%HY�0���xLp�n��̰���Έ���ȭ��CmF��q"�R*pp��p��`�r�Ή���*@K�?��[�����fk��r�����1Y�^�.�+�)�A���g��J����܀�+{�!��r[�?O"���mg�cL�Z�d{EW_�`�{�Y�͝�z��,-��wgd�D�!�o��9�I�9kOV���?��C�h�G��}�Az��QDK���]O�h0 }�S�Jc�V~;�!I�]�y  ��_��ʼ����@�����7���(`�Q��ɭ��PDa	c���Q�"��c-Wi����k�s�b�ؘ7�Ŧ�W^U/���qM�	�2$���9/��v%}7�����<��N���)#5��;��,��o���-�����~2#��I��c���"-�MNp{9���k�ZG&�3瘩�Up��؊�F �.�o��U�ŵ8º�,�*�|�ڱ���a-_��t|3_�ð�J%���%�����7_�J%�ta|[3~�h+;O�9YmVl�w��|������H�P!�oF��9J ]ٷ?��vU8?��'����Z��N!I�e*,�e4 B���ʤ��|��g!�6�t��=�RO'E���z�w�:6�B�b����@�Fg��tmR������u7����P��[t"W	q�u%݄PCNd�8O~.���d�I�Qb4û��b7^��&��t<4��24��Id�]I���<�;�&�l~5<�G�Xj��{�f��QLV�(�C�me�_�۩�و�ȯ_p�[X�Y����y�K��A�P�;�����%وhwu�Ne%:�[n�����A|�B��`���{�?���y�T�`[@*�j5�]�w��������`��Q猹�����ob�,jEW�hL��ĠoԨj/��Őj硎���j�4]�T��Ydv�z�E*CLaZan�Z��<;I�*]�%hL���;F��|�"l�����BK{{�Ո�8�hȟt�iQ���\��k�'}����R������̏1�R��5c�#3����C�{�GZNX߫A��y�Yĝ��*�µ��҇\)��{F'S;��Ck�GE\�e)ӵM����!IT�Ӆ1��̺c���3�m�y��
�<xk��P�~��?
�̜aV?�'f���Z
�1��7�Eg��('dr�g�&�p���`���/%�J���C.�	�5���D-L޵�op�?�EC�͕E��[��t��m'�7�T4�u���)����'�d&�Wv�ں�ԮP�zĕ.R`X��V��-~�d�C����3EbWi$C8(:O�5~��O�K-�p͏�J���f��]/{�
ʶ�h`�(����"~V<C�]A�cre��Te��"-���
�G,��̸H�2�m�z��P�<���DLT��W�nZ+�%�(�IP�%�FA�aH� ��V(�T�:�#QS-9����B��s��5����z<����4�@j���lL����-��8N��L҃*jȎ�$ *��3I�ɃW�ޠ>'u_;<�!�K�I�j�.�>E{"����Wp��u�ցR�Kqw� ��;w���R܋C�(�N��� ����\z����1���kMYk?9<�G��i��)i�3�m%_�l�������g༈*Q�[��³�O)��R/B�&���3;��`|?W`�>��>~���ō��L���oܞ�+��N1�D��[i������8�S��x[f�Xc�i���W�͗��`�G>���Rj�QJ����.�^�<`'�����Kj�r�|'&������5m$DA y^�x+2�J�ʚ�(�5�r#�� s��P��R�b�WGܽ�a�����ߪB��Bu�R+��o��
TZm|�eC2���l�T<�r�b�xlU��-�����&�b�����R�b�ҔF���}�~�k0���`���0����l�-�}�>��l{4�*M	D�i������nUx\
߲�\�=I'e��A2}�{�a���@وlˏH���f��e�$*1����A���܃�[��zi��,��3�Hލ$��X�ܯ"�鿯�)�/a�|��rH���,Ɓ�?��K�k��יO:�?r�-���L+�NGݚ���W���,"��1&�	ω�O�q�ZPM�`g�R����3yV�E�la�O�T���I�a��6�ҟ��e�ߦ4�>�	~�/O���l>T~j��D*�C��T�5�4��V�Z��;��|�>IY�;�q���Ç|î��ϜC���WI�i���x����J�}���i|�{�V�T]��'C���s���l��+�<�Wd
��<��=�%Τ6>b�酁)���g�C��Ul�JC!n�$([	x|sh:!��j!}	v��"g�T�΅�i�B̍O�2ظ��]�M铘��EX�'dڂ��!�ʣ���l�g�m�1&����^p�M��#���v5;јfڠ�tR��a�'��u�ģ--5�U��_�]�,m��<SZ��"�vx
��uj5�qWM[�f�c�zt��\ۭR���/�c�3wN�_4 �u��ōo��_S^`/{^�4mUb�y��.��Y���d��ڙv�<���e�e+��f�M���
�2O$j��/�_,�����q�N3�N6�?��/o��+RO�d)Er�y����2���_���3���gv�+;��y�����]y��	ח���6f|��j6�$�o��K�Dt̜,=��Y[�+��K�IG���J�rJ�w�(z�c�b�\���Sۍul�J���R,����ns�ӻr\#���jP�6"��|��}���&���veYY �6�!B��I���ڻ	��f��3[��kR�W������ɖ��D�㘈<2f�1�c~�6֩%�ݺ̜_N�ƻ�s�lE_���Y������:�T���m���.s�ki�m��U��� ��v�*��3�r��>c�D|:��� հ³)Kuѷ,�4h�5�/�L>{
wC�����ޣe���D<�ށCG�S��9������o]���:�ƙ��MPS�%�ca�{z
�x��*����3o����
���[&��!��	K
�MCH��rK���@iu?=������ۿ�-t��L�+��F��Աz�՛�����A�wG�ʳ����k�E��ޔX��R�����Tx"O�s�����O�6T���8���vaOU���0t{��I8N�	�g��6셔�����y��|P�ۢ�j�zQ��f4O��rlh�v��ʃ-�����嫧魊�{Ζ��b�K�����/e��&��v*���;�6S�Y��7jk.ϸ]2�x�I�?7)~�I;#!y	rx@�|*�?~���Tc��
,��F9���/	�c,+T�uW���B��l��U�����k�Z&��TtN �^Ó���E;'ص�z�r68��,4�	�R�x��x&&x�0|;h1���/���w��1��bH�P��o�x����̋#"�db�Y����>�V;��c��>���W�ţk�Ä9}����ƣulC�}����Փy�$��Y����^wVFc�bHt��F��󦂌����f����^�\�$e��G/P�Oid�H�9Z��ڙ�'H `����"e7`���'�
��
/}����e���8�^f���br��e�?�������2y]c��x�PS�7>�Pi(�W%,�PG����R��.�lq����D�	�}5.K�� C��=c��>��ll �t)ܙ�`�k�`���	�U�B����I�y���)v�G���v�ǝ:vV�M��H�ú��!  xU�������
˙����Ej�"&���n=�RR�zLMmѷ9�<�P�PV��
*�8��B#c�\Z^�>o�Uޗ�J<g%x*|��P.&��:��=n�V�v���S��%o��o�7��٧*��С����!n99�a�t�,76-�&�o0�R��l���&d���|�T���������N�Xﱭ�{c��9���A��؃�k��ʙ���X�j�Izoc�^s5$�V0f�׋���:�+��sޢ��X�e�[#w�m(Lv��Z�|�}�/�Da�'9�a���ѭ�ˀˌ�Kd�H@�ޡk
��,)�t�J;�O�#$��%�<�8DJTk��Y�����#�:���Պ`���5Cս9��V�稔])l.�����=x�6��%v�Kְ�8��۟q�7�b6EX�p�|s�� K���ߣd�qOJ��_�Bd��_�����C�u�X�/2V�|�V?n�r��;P�]�Q�TVI3��-���)�o�+����o`� �.�����f3�y!��3�XBқ�W]�]���i�����_���/эB�qY�~����[�dڠҎ�A�9���tK��hls�������������?�ō������!���*��y\�C����q���=,�����66B����M��$��7��:��9MOf��JV^n5�R����æ���MX�A�v�#ں��k6�z�/�f�bZ#���AU���)L�j��s~b�)����v�z��x�Y�h�������&�ٱ�;u�����$�'	;�-�-�n��Ɖ����
Y�Z��׍#�u���}ɇ��Ly��ɱ�@���M���̋��YCk�qca��������qQ��
r��D�x�CY�%�V�_.��[5
�Z��<eB!����O4�g�����Ű�� ���
]�x�Fs~��u~��)��B�-f��Ձ�ƿ
q�?0��7��MW�����'�x�'�کň�.���Z^=�d@�_�>#1ԉq���%+�� o�1���n�S��`&^4��A���G��w�J
�>s�CWn��ԁ���σ��b���(��a�uNf��R�s�[�-��،Mѥ^0%�%�8Ǔ�\��ϻ�<Zˁj�~�c{��Nes�N��ϲ6�n٘���ZV��&����E�Qnb�N�&�ao[�ӂ�+@����*�l��E f;���Fz�	���@>ĲI��Wؔե5��f�3����	����1�ê���ʛL:L�2"��r���
\�K�3י^�^$XU�,���Ef�z�'�Ҩ�A��~&g�5Z���i��QI,�ߩJB�O������1F-�Y���}��w�l5[
����p$�M@{�p�&(-���[_�Z�:##\�SV.َr�?اfӴ5C#,�磴��ԛ0��ͱ?v���D$<��nost��RO% jSA������dy���>ȝv�*+)�(®��.r4|�2I�󧘈z���	����2���Ջ���A�U"l'���"���~ǐ���,�d��SA�:
���\sl�Q�`�D�����)��Lv9|W�p/���>���h6o�����,P^������4O5;���l�{�߰%��bm�sW/W�ה����y������]ZU8S��	�g;��) �=���[���1�df���XI��A�X�y��[������>����2ݛ��S�6	�pB������D>�Z�I,�5�~��L�F�#�xш{�^��"�k���z��.6�a�������!�1Tռ�(��y�b:�-k���E�4e_#r��;��-�r"jM8�Hۑ~?)�@����}=F��g�p�y])�-��ɼ���''8$=��W�cDC�Ѕ�2�۽�m�&&��w��-LPC�a�d���O�&���1W���ʝ2P�VoK�Z.�\��"���!�Co0D(�Q�o��� �)~��H�b-,��U���9؃lK�V��}�/I�b�4j`�jL:��Gnt�E	��Mߊ��mA�K�K�+�2����&����CJ�s��w[����[Q-ȂB�.Qi;?��Z�(���sJ�F��KR�̏{d�}V�����#�y٥#x��n�q�,�hzC���xn=Jc|1a�AR}�Nߴȍ�zv�O�6���>���.�7J�@c'��N��>w&x���[�7�\��GQÒ��|�zĂ�/�c��\N������Xu���7�����T����!� �}�N�'�r�g�W�z�.=��d��D�(}m�Zh�x�k��>e<=0�5��U�uIZ,������:������Ki��S���I�Ȋ`Y��p�~��%�.^?����T��]�,�����[�G�Fw&���j�5Dng��S��J���V�����+�5�i.��!̂Ѡ��V Z�yO����j�Q��pZV��(+1�g�|�+�OϑM�N&�5�/�w�;/�s�c )�t�6��'���O��ח
��ٮ�%O�?�τ$��J"�㦅�BQ��;�`q� �0oEU_��YM�z%�#�s�o�-^�@f���v�6?;���IަGJ�iG���Mo��Tu���r	��ݝ�v��ְNK�O��,�Cm	^n=��D
~�<����w�W���\Dtp�6¨��r�i[�{9�*��z�eaf9�=:�c���t�WR岞��[P��z��
WIzqi��#���C�̥I
����|6Œ1�(��!�ޭ۵������W�C�����Կ�tm�?��j����Nĩ�]�x:9��mO�<>��jS��V����2�T\�nC�TG�`�}+�7ʉ�,�^(��nI����H+�/�	I�����%��0�cȿ�h&�M�`'����wLUS�ő���ڂ����R�5�]�mk����<�OA{��'�f��e"N���v�(���ͮdT+2+@~���
�k�ժH����;�}��C�;3�_����2����Pa���/DI�N��!��f���43���������DaZ����[��F ���
�?8[��/��q�|j�V�^���X(��r�S����K�$��r�`�dVL#�!�0���2�DFKO_��0��/�a�x�X���R�f�m�/�_.��f*�-���oԳ@1φ�I.53;=3����y���-7\|�pr��+�=+���l���|S.lcƠGa� ��@16V�0C�6	g{���c�8���1��~{d�L�[8����T�fl��O�̈́A2]�Kz�{%$,JMz�p�PW䉴<�5님������;ZO��	�p��rx�/21�F�=�9��t�e�yr�h���yO���}��V��>c仞�-,;�7NhEO<+�fUyU����i�͢�ߙ�6^��jΦB�~�z�O5�:�k�m��̴�e��5"��ѐH0n�4�Z������[��σ'`��(1�ɟLR�Q��aW��g��g^�F���B�*>��ŦW�
�a�G�z��$Mٝ8v��Z�^�8��6"l<|���Y-ەb<�`�[��\���u6�ny,��TA�W1�Y,�o�w1��>�w�y���"<YL��T������ �J�#�kC��O�n�>!`lqf2m�z�Pb�r�mf��ݒ�x+��5�`PJ����Z����gh�X)ڌuye��ȣ��c���.
�Q���u2�RHV��k�2;ү�lr�A���ɷ�n%��䋿tt*!Ie�6���ws�e������v��j�O!��9�L���"V��K��1~��H��	o�������?�_��2�V��hƛʘF%���J�W��D�1�Y�Y��$��F���x�DP��,[&x&k���׳����_�cօ���H���.��a

@�S)�h゜�A�~範I	Le��� ��a��S���"8������S�Bo␅�@?�����s�:�w?�.*V<����i�6��s{9T��b��wqU���5o�h���q$�v��Х;mV�S���N��:�E�۾�?�x2�=	���Ebڗ ���W7����B��4��n���t� '��(a<�Fz��Z�%�D�z��o�x��@O��ZU����gļ�tw�E��v�^�>2����	ARcU�G0�n�p-dcPz��M)��g�c����	�wG.j��f���.F�o�Fb.$11l�$-��f�$12�H�:�f0�	K����ޝY?8��P�X��ԌZٶ#�U����;l�mC�z��I�݉[��|��J�d��qK��p��%(J���p�S���/'��#�3)7����֥������v�^o�TqhD�����wJ|l|�6����qUS�Cݦ�3a���>��J��|hm��c���Da��u�/�<�zk��Sf�]�I�պ,����;B�욌�R��E�1�-�� ������h�}��Ej�����H+8dmow��-�$rs����!� �mA$:�`�0+Z؋[�|��� �H[�ئƚD�Kg:�>�
O��-�n��(�Ѓ;d�7��*�����~��r�^�"9Ɵ �w��G�4�� �G��&�:w�:="��c�<@s�5�/�o�ot"��7��c:�r���X�oW�����hf)�?�P������yJ�L�@�q<Y��m��R�����6,�r��1Շ����?�Q��6�4�f[(��u�lhR�����`y�h��(;�=��b,
�.v�u>]�a��t��ٝò�|�hN��s��n��Ds��%�ێ�(�\B{f~��wP�;O]�q�e:��|:��ñaX�<�jfJ�!�ߪʝ�&�#�~q�QA���nT͝�ݻt�7$���(��3��꥖��GM?
��@QR�_�2��g17�͑aR�SB��0�"S�r��_��oP8-�p�u�{K���^�_��䕄M~MCCH�$8f�]c���n�;yɑB��{���.�����b\�Y{c��`h���	���<['��t������V[h�����Fhpu�AҾ�O,��������Xt��K��O���1D
*���6@q��^9{W��xd�`�B��5�fݬ����D�N)�$:�,,j:�����C���w-2|K�J	�(��yA!���WS��NV+l�5 �$H��'�(�c���_L�~��~�JF~�����m"x�vw�������(2qW���F�U��8b�+80^e̼�Z��c�c��J{�$҃o���[82�y6�8��\�f)�ѝ�恎�wK���=������^�형�ƚ���}8z{Qw�阀��A�|��nj��O^�b��[��l����i����#�@uAS��v�lk܍ƌ��RY�iS%�@����7�:�nH�jxO�q"3	�h�-r��h� �H'گ��=�C��o�H���^57cb��p��(��Fٻ`꿃G����_W�(M��~�U����2ic�ǖҖ�}|�+��E�~��[7�?��Ǻ�����a������!�)���w��}�����m�����!G֯�>�v%}�|�H���A���Ͽ�+�S�X�M�/���H,7;�p��.D�G���=��q�W|u_�L �r=1
?�b�-s��8?�;�k"Ra��D�)~�F�F��N26+���=�K�6Y��E�w��+����k�D\9���N���`?|l�k����)�����O����S�:RUO�=�N�]K�0�����@Y��y!�J쵱��������%�ٍ�9WA�*x���R�����R��[6νmϨ�K�� ���m>��w��˧p0��t��4t����tۭ*(�͢����O��� վjs� \���lP8]�!]�c	/4���j��X�6V�7�YYPOC�b6�M���b��h��. $}B^@!�Kv�g�d�X~���`�}q��!���z�NE&紦�ad Ҍ�z�Rd�Щ�������3�%�Y��\�>�4�z��NP��D�-�x���$���ͿZ5*� k$����b^Tբݔ�P^�x+�nt�߄>$��g�k��0.��q^�.�Xi����)��VQ��3ܩmV��"�)�D;���3�O�/z T�ن9�5{Ĩ0�V�M��C7�ZA4x���T���Gh���2feb�or
�p����G��|�Y��j[&8K���_1��	�RG����\*7�+b����e~4yqud�HZ4������a��$���=R��֧���l��*�6٤Q�#���e��Y��~�-��Emn�I��'!摾%*V��w���	�4F�Ҹn��r���	D�o1~��PeB�?.H� �<3����h��?�Gy���K~�����u��'�U�n����'+�[���c^�k[7U����Ǜ�>�BH�Q��b(�~ +����k��y�t�[=�.�Coˣ�t]�"��F}@NF=����T�� d�9f7������4���ףb��'9�Qt�8:RgE���KEUn����lϫ���=JkH L��7��d���>��)�t�y�<~����e��R���曾ֆ�3��&�,�_]W����	m��%=/}!�aZ_�s�~�xs�
I���gj!�5�+���<��Y�<i1���=�Q9K��"gD�6�mS�%Rh��q�ӧV�@�-�^�w�"Z����G?��<�j� Y_71^�1� lM��]R��I�+��/V�#Q�١�YB�����_�ں����<k���ũ�11=��� �*pO�t�ů��N�?�+Kl��j�>��x��#�qm8�_YQ3�ӻ?�m�,%v�0JN�����B����(����^㆒�>ip6��+o%u����֣��3�]���|j�������&�1]�F0�UϞ�|��I�[刦^�]鑢�fEt�W���e���Rq�^�T�w ���P6�z`�e��N=&��/��5�z�?Y	��j�_~ ��2�W�r�⏱��鵔���G"��a�|���B(��G�})�Vъ�!k�B�M��/�'%i�[tޱ��ݵ��T��;u�/|�y���\��Y��{��0d�%���fL������Vd���m�;H�E������$�q��W�'%�ua����ĥ͎W�Ǚ��~\��o��U�Ͻ�2Г[᪞���~��s�S{�2G#��WGǷ�;��|UY���&D�S�g"���&:/Z`!�(ף�Cn<��{S�J�b�w~�����!�4��:ʱ��!Z�[�ِ�m>����ͫ�A����QL��X�����R��m�^g�s��;��3c�v�C��{O��$�X�H�Ť�f^y-�ϦV�;�E���Z5�2����"��Ī��f뚢|�r���W ��L����6υC�l�"�?��6CN��Hl��[��e�����ٿ�<��xMeR�C�����Fѿ�n�C�:p�����Q�+
��eT,�?�f�&�������O/>.۫��Sc�����a6=s+Z�o;׶�p�b��Ѽ��Mv��`~S�=@*��-�bͷ"� �~m=[sW�g�n|4O�B�����h�1fmQ�P�U�á�L� ���F�]�l��yt����I��yQ�qk!�j�7�Gf�S�]���B��V� 9�b`��x��QH�[�^9�1��gw���%6H�z"���Sf�w�q����o˙>��H���Z�i���<�0��w��<	9���+���,L=����N=>3���2�!���+Mչ1�3� �F����L�~��^:g7YWS[�S�{S��_��oߎ]��^B$v ={����Y�gz®���ql"?vz�	U��"��.��K�2D�E'�'~+.�Z9���gט�wI��D{�v�L�QM� G�viŅoh�����k�S��֝]�8	OAWܖ_7��Ki����6i��5��Cb��-Ò����s��Y"}�pT�6O_ U�.`E�K*/y��^8���/0��y�L؍�)E����~gI����T�ޝ|=�mM?��X �<�]�����+>����Σ�8�mDMs��$�n^�����"t����o�6�v0��9�o���r_�17�����گ�QwG9��-
�:M����a���chGM�m�Φa ����⺃r,3���^zH��?ߠF�]��ax�j�s�2^C`d��u݆~A#}�{��V�Di��}@ �D����s��uފV��@����,~���r�l��*)��������T!ƅK�7:�o��nq��i�����,�P����}�!��\\X����R"��Wg�R#!1}X��������@6|A��d�ݬ�����{�b�M;Ь�h�n�tϤm�=��ӛ���Q/�5۾P�0��_T��P����5�.��J����b���xt>MM���6�-	��i����?����qT�(���3�渊.7�:�5���eo|��f\vMq�i�:�3��vz���Q��Tz5ch�/�0�t��7$��Q��������g�+r>"Y��8��Te.%;�7�
��߉���ڮ����؊��׼��쯺`R2�U_�3��O]�:?����*����/��HS�h�'6luf�P�	�@�Md�I�t��\��WZ/Z1#<0�]�_�6�P�j�J�Br�����كP#����is�#�I%��sD��1\���U����� ��SS={�_C�3�J�7���	0>�L�e)�U�j�b9�?���]��"4�顃Kv#'�4а�wl	�aO�J�L,�<�E�u�n���޽-�����Yq�&"(a��t�8��n]�'h�����0	��٣*�Me�j��]�(kEP�/o�F�6�t�(��<Y:���EWv�ޤ����t��$;pӦW���x\�'\	r�&���nN���w%�{wG�S��v\)f����x?;p�e瀲;�.%�f����t:�@x�q�r�:�a=6���2x��v�%*���ʎ!e�]�tM׼yn��.y��)�M\"7�rC4�-
�v��筥�C�V@�ge����X�m~�D��;�m��bG���`6��A����Ҫ�zO��̛��P��.^h��<�Y�_c�Ux�d��3�?��j����b�Mf�h�)��W�v���>4f�S�z�6M���֢��i�̔�7�vj�#_��կ�_
}�4 ������\�~���#����5��ýz��p�!��u��Vo|����[�h��Kb���^�̡.l(�`f���t���O�x9]K�^}��h�B8{���95��nߛ�߇���\��Ů_����A�'s}Ju����X{�qtF�����jUh�r�;6�o�	E�ڤD��#[/7�\��r6��ϻ��<�9�(��i��-'�!�x��L��S�h�!.���6u���N��3*-�X�O�]Hz�������KX��Rb	g���i������z��#�Wm�k�;��-��0 �L�������z"�|�}�ɀx4��Fu�5'��ʋ���MҤ�Y��љ������6f���|YF��A�[7�щ�#ӑ���^�����9o^�6E��zA"�D�U3�;�f���ؚ�T#�c.Uמ%K����VʀAH�J��^D�X�!�����mK��d��G��ݜ��`�$���\T�ǅ�N�o?��j57]z\{������j�8�$�� ײV9��Ѫj���@z�ht�����ݬ�Ӄ���һ�n�-{)�w����������5��Vܧ���0�&�f��Ԥ:�I�Z�Ë�3b��8x<E9+E!Q�[=���1فl�+�20Ə��7�Z����[�tϛ/n�8���X���Пl�S���6��Ӳ M	�H/:���z|��PB�aMb&���
��v�δMK_�h�nkJZ����6��� )���]hד�Ǝv y�K�*Bq�l��mRT�!s$i)�M����e��Y}~[�H*ߠÏ��d ��ޏr�7y�6
rO�"�F����2���,�����C�n�v�� X�U�ڞ%V����A(�*�=z��"����(%�rx�_)�������lNU2�f����WBd�'�r5�x����@�b�6��4q����o�4�R���������>]o����+$H�r��?oH���ϡvPK�5o/�S�=��u�[�Mf[�R�/p��)�v�@"�|7�**�#�B��8ţ�wh���ՙ��]�G�����(��]t)�I���ln��+�;mS ]6a����5��]Ҧ��ͣT,E�et~ɇ{�/�drW�6�����|hymR��G�\�B?�x4�B�>�2�'L���&~�KҴ��tV��<�J6i��b:��'O�����m8ylA%��<;����J$�����&1��PD�P|��}�&F��F0�E�\w������b�Ae�:��o!Ӥ��-��h�$F����a��I�����K�^p��� �b�\�r�O��6z���g�&�K6���<����q�m�ǽ4�Y�ލ��M�]�.��\gQ��yֆ�%5�^k�"u��)aS-鵳K��*�ϟ	���r�{�e�>BL��k����E9���6�^o����Ҟ���yb���Qe��A]���*'���i�0=�@���R��	{���G݃�����j8*�^��������{&��%�6_�\��n+�Y���9�򺯒g������eo�>�*����f(��`i�<k�AΜ����Q~o[�0��=���ۧ�<u�n��m��~��#Y�PWL�nD��7�}p%����j���ȇ������s�_�"i�fr<��[��Zty<^��~Pd6�ߴ�h��2{�ȏ����Q
!����GO���E�h:m��S��V\�d�n�i9Ϙ�������맘�~�z ��Օ��A&@�`J�	UϘ{�B;U7�ڬ����K"ot�m�rtm�&m �g)�3si�[ep{��%��:���6�ݠ��'Ꭰ\8d����;�������6��df�V�섩�c59Y(��,�8�Z�н#��ӧ�2�1� ��l���gl2�����A�s2����嚤kX�Y����0�:=?Kc5��2��T<��{!f���{�'��ޕ�����}BtR�{\a�w^����&��W����%B���^u�͓���8��i�;
�U�	���8�p0�`�d�Ɇ�}c��$v��"��I�p�:�]��<RE��j�u%�f�%h���Q�]t�l{;8��q�݉^D�R	��Gw�mB��]�L����jpЛm�O8���K�"���+cp�e-~���ag��W�=��_��	HިȒג2#w8'<����}&�m�連<`�ED:����&sg�">����^���.{�㚚�i��5"V$=B��"����N{����6�W������l����0�H�	��>(��W��b�Ju~6P4N�(,t���w5���w��+!p�cB�L��W��H����nw���=:8���t8˱a��@�l?>ἔ[��zڹɀ�n�L�G�����p�<BNƃ�"ۼ���8~����i���~D,66R��è
�B*��9K$�V}ّ�,�&鯗 :�kK~Q.3f�ӆ%��yK<���e����D�����Ň�\�?�b@;Z����.�[Fw�,�]�^bP6���Cj�,uI�$��o�;1Wv��4�3�S���|�k�5z�A�>U�Uiē7&�a<�����#v?/�q�G����7��xwO�n�[�M��ٴ��>�=o����2�ل�E2��u��W�U;��U�.G%��� ����i0��	IWVK2��Q�Ń�/��N�op��EPVŕ�̻�1�D��x	�lyg�$"yC�&u�K����������p_=�l|�@kA��!���p�D�t)]�)�Kv���̆Y��R���a��NZ2�Ê;��G���G{��k1���<ˉޓ";�� \J�߬�=�7�Nx�����2H���<)���=^����ϖ������O�S\�fU�:��L	G�e���#���{���\a��8W&�g���L������U�e|]7|�8 �$����[ڲ���D(&Rw��t��FN��f����v�ʗ�}����M�6��.�?�.��1���'��^�O�$N�"\�v����(�dpCO�ԯ���6�{�L�X$��W=@
G6��oRw/W�~���`�y;2�>h�h&+��0�l���RWJ;�R��X��`�04p}O�? 0l��S��Dߔ]K��n�k�b�\,ŝ�m�N����w���6�"�0#�$ٖY��1D�
Ǚ�V�0�?2R��04�����S�O�>��.�n�FsT B��33���.W�t{�[N^]�d�RF�|��\�:n_�]i�L7�Z�ٶ�Sl�*�w��hvPʇ�<��|7��s�\�?d�0������{��@�{aYsp�ba��.b�tr�C�+��"��~C3ÞnK3L�eo�b��pd�1��l�2;���T�����CI��/E�_�	tsF��8+�j�e%�}��ƃ�>��M_Q�y%�Ǿ�l2U���Rw��*rpjӻ��4�b�B$LS� &\�՟����N���}����f�jr�%��-Y-�{�c�Ę֮+��L�XCTi~ګ��+��_��9va��W\��G�A1�l�
N*�2_N&�:��#���w�����/�_���]��*W�E�h5�K�`��:���j�m�����dc�s̗�0+c�[�����]��ʥ��B@��|��m5��bp��A�F�K������~[�� ��N�K�d*�Ae:��ڠ�Z��l*��}�v����R5Zs�\a��]�v�K2����|�³!1���L�!���F]-7e��0��1-;�./���I��׉�T ?��]틕�7,>�d��4������9����Hv/m�h�%.x8oct |Z�%/�H(�-Oށ��D�:֝����.ZW��
.Mo��=�n�M�,d$��nwb_X"|
��:��=�����X`BhQy8	m��.�D*l��ˠ6Uc��I����uQ�m��+��M�|]x��!�cj�/E������AHR��6��������ແA�(s�NŐ T�s��U�]����^�i��4����m'��w��OV���A#���K�f�'T`���m�!��1��5-�<CY狤���)���W毿%����R7h�ViH�Hd�������L)Ju�D{���R MI`g5]��\A7�?����o�s���v��<�~_�[<��qи���_Nr+��;w ��߶u	%����ѴTZ�_�p�n`�Y�-�N�ն�{���dz��н,�d͐V��D�O�4��R�eU_� �����1�b���U�Eۤ	�!9�% }�������a��o��]��i�i^Z������Ǆ�yK�����P	�g�Y"C�{9d��^�GG8E!E��]�|,��Θ�$���ܒ@(A�N��y��X����QX8l2�?Qӿ���%bܳ�_9xqK��$������q�~��,���VʃU:���vnޱ�2�����Ӎ�y�q�g�*$ӽG���.�${F"nsO�"�D�_��$.A�/\w8p��!�\��A��
�1T J��m��	i�zτ��_�jG�}ݗ�|���-��Y������w-�;�.�g
y��S����a��HE�4~���_x�Y:e,_�"�د�c����Yf�ļ�m��inY�|T�m�����"�S\�;.��uŮ���zy�g��$���n��%���ʱ�}�z�-9����� ���Vk�kܔ��Gr=�?�)��-�pP�e$�����R�O�%j��(|��ޣY�@E�F�Ry;�Z]5�5p1�y�-����j�4n�v�?o��[�Xf�t;>������]��=u(���!�] ��ޮf�"��?��ծH�2kI-6[(�t�urNӺ)D�����v9�b0vLU��X��N9�T�;�@/��5Ț��G�����f7���29˿BD�ՀГ��6����I��n�U8l�x�6��Ye�ƬَE��w�G���\�>�%I�ߕ|�����e���5
;�<�����^j�ﳒr�៙�pڼ��.?ZB\H��5�,�I���)�u�J��l��6���ɽfR���r�Zb�� ��2V�)�΢�ͤj�Z濦�V�|�Ii�����y�2H�am~9ГT��j����:*�FJ�n6�9���P��[���O����
����� �#]�H)H	�-͐*��1�9 54#���9t� ~x�����9`����}��*SO���gYcU�w�$ݗí����gՆF�$K�)�eO��=�ϳ�+4TNPF��e�;�h�v�<'��(̳��|���e/�H�yJ�=?�牄Ξ͊s����fp[��(�\}�gWXK�y.�+UC����u���P��q�=b�ߣϴfH-�>#kni/o��"�!��$��g�+C�])��E�*��չ�T�R�K�������|�������h���[���r���b^��;��H�3+�e�a5K	���M�]�����K�'l�Nl�E�L�6>����.���֐����ШǾ@�C��'g�;F��u�^�i��+��
T 
m�WQ��SR��v��lB�2�=ШoP{�]5�]s�V��V�FW&mz;�<�Jް�կk�wG�p�ˑ�������α1�^���� cĩ_g'���l|�!��/�k���I�{K��Zv0�[��|Ǿ�;�FYV�|�E�� �⮒��N/s�2�]��6r�173e�b�̭&%6��:�
~r��b{T����ݢP����y��52Oڭ"�ʆSz�t�R�V u�w�yS\���*����nT�C�B��Dς��ԃ�L�k�Ȋ*���0/�䱧��]��>��_-�������?�u��"䐤%h�r��L雷r��;s�$E�ݍI�)P���,u���������o��M�)	��*NÆ[�)�/ַv�r����]�[�/�$x߇�N����<���h�hS�Ǘ"���41�|R�7������&P�/�a�g�z����7��_VF:����j�ƥ�i/�W`�+�r9���?�����_l<� �dR���Y��ȕ�`�v=U��=��/��:�S����9��Qbrja�ݠ����<ǢX�e���Z{o�Jo%�G�I�ͯ�Ԥ�ά�x�j��b&ƻ���|�a�y�Q�5 �_N�S��>w��L?9� �K�;�$���h����pI���?C����:�QA��N�ǿ����]�y�7�M���O-ɜ�w�&d�
��%5�x	�+��.b_�ZC�.�u����ʕ��
���gG{ڗGY�=����g-t���'���������+Eͺ/7)��/�MHt���c;*�!��t�ˮ�zmO?�f�����13?q%��Q�X��`��,�rY\��)h�}2���F�}:Y�Rݥ�gg��g�ۨ#`Peτ(brD.S,����w���1��܏��ؤ��ہdM�NGk��l�P9�Խ���-�ja���Y7s��6��e��V�G�v�����x�Uc�nDc���;���+j�E�U+Ͻ^�ˍ��7����'���L�qX�.��|r��1@�e��o(~���	�ߓQq@�ʈ.�L�5�p�~��,�3o��´�.���T��ଭ�X(C�Ң��[�¯�.�ݴ�;j3U&	�q
H�|���ڧH������veЭ���"��
�_7��̲&_^
 eK��F�OW}H0�[����2ۦ�%���!}�A\u3Z���Lb���B��-�z7���Iu�WJR�	���ax�
q��z�8q�~7TO�)��3s�84�X�ҫ�8�\y-^c��˯*n���l5Hn�&Ȗ\;Q���G%kl-�tG�&,���1�1����ͼĘE �`�ڼ &�4��M��)����Pk&�E�󜃦��=p����rϼNh�����9���!#���dE����$����V����X��;��_�]Јx(�\_O~I֋�qZ�]�L��*���X�R�~l\�(R�H�B!�d�)Q/�����cJŮ��k��q�z*�fN�IM�*�Ӣ����8\�l�lbz���X�����0��?J��u�&����E��=�L6
�|Q��'$9A�:P<�,1���/���7!��OZ&�-�΂�`�Z����<��ɚC�|�`�=/v��M޵�JHc�Y%9�Y� ������3Y�1��!)�#�h9���
�{�*,H:g�A���u	���ZY�g`��Ok�\��c�>�N��g5�Ѳ �0�.��s[��rW���"]��W�3����e���X񙮺"��CrIL{8�>q���[�P����k�߿l���K��+D����]T]	�eSm��g��J�u���`�1��I8��,y���T&Up���I�	�hm�G�^��Wfĝ`�JIe%��ð��X�}RBC5�x�D���=ӻ��}��<P�Y^����p-�W�f���3�����jJnv  ��f��h{���y���מ����<n����,(;���G���ۥ�O��ݩqIw)�=�NY%��c;�؋L{���Ky���f�� �5El=�9dR�B�&�A5rŀ�3غ^�۽~@a�ݻ��`�"s������xԌ;*��~�4@�)�G4�`�{�nC��M����'�2��0 XX��i����/4��c*�ڳi:A�,��f�ޖ����:��=\���D�ގ�w�kN^�x=��qq�1(���W��ѓ�V�4���y�s0�e�W�a�S���Xx+�y0uK�uu��w%�v�wӉ�Q߈�l�2׃;�?��+�8St��-����|��GTf�_�.�B}}y8E�طEm�U=�D8��2k��|/%6�{N�FM,ڱ�<a?&�24w�ٴ�������&��|4���8<��掕���
8|����K�8�;�.������!_wMm�&��c]0(3�(��y{�Ҵ�PPJ�.���Ş�F&�ր��<\X�R���Lbd��L�C*��/��\?������k$���Y�VHϿ�4Y�o$u�F��a��Dr�z]�2���*$�6+�UU[���_�B��U��9Lo��D'���_n9���[1Ðg1�� ���W�{e.m�+�����W�J���4c����O*0� 4�y�=���!�Xz����9��'Q��#�Z]W�ʏ�|�% (�Z=O�&f5k�����vO�_v�tZi(x뤫�_i�����9E=W��r8$���\ďg�ب�u�h���8��\�bS;��������&z_�����������l����ԯ�L�v�L?
�FUu]v�P���͒S�Q���(ǿQ!K�<�����g:|�ܓ(��F������ &��}꾘�	YD������X1�����p?�R��y�9��&�����'P����A����lۯܡZĚ$6%H�ƾ�<�nrn�Wӯ��la/�u��ݜQӄ����6��3ҎG֜�n��mԟ������ݣv+e�BvV��!��6�ė&)о��D'�S��AŌ��(�V�b�U�1P�(~p(IG:]�Qc��v����Y9���b���?�
e�﹯�
��	X#IQH����nVpx3��L�ԉ㺊��w���$�Z|* ���򭥒+4��d���I�ؙ�ȥ��M�Ji M�r����.��Gk=�q�ȕ�MN@�5��Tu~�I�+�e�SK�"���)6�*�P��Y���3�;J_�/$ A���j�H
s��Re���eV��F��F8A�q���yغ��ȵ,�#ŉ&Z���V�������h3�4��R'�v�Ϥ1zVޅ�0A����~�<$Ic�y�[���f�@��x6�8�|n�#�(�$`�f����\t��w�{/,�(���mE��bUXL�:W 򸴻J�+Sg�YH9Ʋdw�N���]M}������2L0E�^�;�
Y};�}�`d��Fl0�9K�x��,��L�gz�m,���nJb�F��]��)��{�B&��7
��+��k��.�x_��,���$^�5����@�����_m���/�t�)�?�U��iہ��U�L����$%�����
0)�
匹�=�؉��țٗ�su�)�˥ֹP���?*G���[���fzaԄ�4�BN���q��cp����=���|��%�e�Y(��"��M���s�ˊ�&.�#\�}ܻ � (�6�-z��;$2��������i�%���'�Y����|��f����n7��v3�����Vx��e��3��pӵ��_0��3,|��}?lg�z�>n�5��~z(~�����N�Z�q)��\r�\?vim��a�lN��E�H��Vn�܄;��:s���Y�֗{b?�\��z�q��<,KĭC�-��p�9{i�f�%y�<��ǡ;��]q.�1�[�M�q8\+-��7�p����ܴ�z�����(�`{�*,gx�
b}��|H�^�s�h�����I�z4<�}��f�8�ޞu���_6�Z8 ~�/DWY�W�[�Z/�ʥOJv�w���,$R|�K� �C����fe%EK^ָ%��؊5F�b �����qA�cARIH��eR >���-V�樏������</c�����u>��J
�>�v[C�_c�y��m�����L���Lo�;96�U�ҝ�@
���ϵ�!�hy�ÑϹv��gK>�>ы���vi3�*fX�m�Ng�А���xmj'�z�t�?_�ΞQt��7�w�������m=C^7��o�M:�@h!��^�བ�L-7�'��J딫����~K�
��*3�F%!Jٟ+<b_�$�ₐ�C��N n�i�����If��{���|��8T�&` ��k���M��er�U�;T���$��v��U-���c�Ǌ`��Y��|�ǦС��{��x�?���,��Q�MP��2�'?-�܏S�7nڶӨy����N�u�quoxe���XF;��!��������3,���W٢pܩT�tj9�E����gc(����QX-Fe��dm#D�#pҦC��,��>�l{EN=ն�P�ym۟�/�I\��Zzd�è�:Pw�U�{�ST*O����B@s��)�%+��CG��hy?~Y�-�K�v��~P��S�yϻ� ��y����M���y����빅�G���o^h��J�^ fn>�҈wh�.�}k�2����rQ�w9Cd.�=��e
i��#:�Τ���Y�'�Ӟ��>~2=սt��y�l�QWt��R@p��#��=_5�_O�F����^]�p�S��t�d�]���D������]��g���K�˝v���7�zx����X�w�.���U�L?)%�\|L����l�Y(�79��ž�սSq貄��6�F N���c��&��h&UD��r�s���W��6���ݾ�%�Л"�o���(�(�}�e=,U|r����b<�Q7 _�u���>l���B�	�;j3l�|"��@I��������l8r��<���_��E.����H����E�57u	<䀃.xe�*8IaG��G��߹�IR�u7�E��Nq�K��m�d(����P�b���滋�U -�9})�Ϯw��+w���z-��zQv���"0�U�]����*O�/���������9�Bb�^�h29���6׀^3&cD�tZ��?����NA.�%j=��&8�f�՞��̀8Fx8��n�$����o��{c��<e$Io���\+��-R_F��7���R��R��Ey�mR,��2�:]a�9^D��<T	~"��ƻ�Q���Vύ6��1������ڊ�S��z��e�]�N�D�usS�{�mz~����fҗ�-Q�d��7�-��&8�^��wB����$gI��5�[֧�&7��K��RnΑ�G���#�y���Ɂ8��D����Y�/z*���5� ����
�x�7�r��L���Z��r��"vXj�NЙ�Ij�*�'V0p�=7B��:������k�wg�����x�M=?�{���굆��H,Q��E/�F�W���@��N�SvjLGߥiʶ9���8���Z��(���c7��T�zU��gk�u�</�O�����&�(�k4���:i�IR��MM��xy����q#Jk�:����ɟRr㹁��*<Wb�b��@���M�j*��*~q���}�}��se�dY5��k銍<Q�םwr4���}��(�,��@ܓ�=�K�H9-`Ok��@T_������IUۦ�%����N�e��(���{��~{�_x b����p��f�P���F W�%��	�q�U' �UI/'��}�Y�ѓ�&���&qB�ii�����0`2
��% YDocc"ܭ���h�c=��6���#���å��4������W�Y�K����1"R� �M��֐��<���s��	.��?؟�:?4�����o�p%69�^yo3�4i���,�����s�m���e�Z�#<5Lv���^/�M����8TF�(��0�!�5WM�����aױ�D��D�׹���`�"4u���>:�v����oI=/�X'�J�D�h��]*�Ρ����g�	c�f�8����-�_�����G�o�-I_s(im`��y\��U�ə^q,�'�p�|{�n>�"
�(8~4��m��<�yd�sp�r��(�6A�ueb��!����U����Ў~��'	�!�T���a%3�����0a^u9��$ҥ�B�ܟ=� Mv�ȷR;�S?�� �JFC*N��6�B����:�-��9�#�	�X���5�()ť$McA��&�Z�b��|�K@��3{1}_^n�s�;��S8�$�/�ܙ��K����!i�>���1ڢ��Bt����&���x
hR �zˉ�����~_]�c�򽾠�ڼكݔ�]���G��4S���vs�����H�-3o��(5�H�c(*�'����8+�^x� ��O��~7�U��:�����n2�:�d��^��GM�=��>��3|g��_ܺ�bp����[s=�Xdr�t��zOZ�P֬�:�R֋����Q,����uW���������Q���#�]���h�T"���Q�_Yb����:��J�p{fQa��@�.����0�����@Y#��n���������y�N����o���kgM{����c]/Z=I�ydO4�R����/5��q 6�L�b���4r��A���t�J�Z]��3����o��f��v�����  �>U�ʆT��� ?�</����|��}s��2'G#_��x���|�ݚ�gd?�^��#Th�2��W[2�d���1��f�c�]hb^?��[M�� �����v��}��E'O�������ǩ'Iu������.�0/�6EL�팝��7���.7(dzY+��.�O����-טzrif*�o�ҍ�C��P��O@��}0��;Eй�w�.e�>���͵�1����>�7�:���ӗ?n?������9����.��D���c��,<���^����X�
J�˿��J�4c�Iг�+�$h,V����/+F#��5�j�%T/r^K���â��@��r���B��t1 4�,0dw��$�.VGؽW"�ksQ#���j���~��sn�_�Nd�4�f~$��r? ��O�m�#����=�b$�W��5<wٮc�I���Vq�R|� GƯ&5�X�X�;B�L�Š�w;W���P���G����0If���� =��n�D<�d����G�/����տ�:!�� 83�M�olx<w�֯�2Հ���y��=rt@��y�_�^u�H��Jm����a����زCR�Jț��z����J���~�ez��ΆH�k(���X�4P�;�/��:�͓	�*�;����Y�(Te��K}���Қ8
�@�8����ea�[`Re9$�D-�VLr�����+Z���Ѝ�?�Q/�b�%w��0�,�^mg.�J'g�O�0�a����e���ة��ϭ)pF��S�&&���T�Σ��sY3��1g��J��g���?Eu��B��3_���3�j�؅��54ׂ�P�t:���.n���E��t�6�;�c��G*��װ/��Yc �87���CM��Y"���}���Mu���<Sf΂��o�0Q�l�*��Ֆ��d�������%�ۀ�!���j\�=1�䗋��U��[�`�IfM��VVD�⡰xv"�v�8��zi���^�!mB��mtqj��W��r����/����%ޕAxZ���f:�p"���Xz�M8��Ld�xz2�:ņ�v��
"|{�3��q��|����(��d���2Q��Dh޸5ڿ�	=04�,�Rj��/�s�Y+MU3z����~=z�$���Ȑ|�<Q�j06%A���U�b�Nm�lS�t�(ea�����)2k�$�A�HM�ͫ�1�{�$��A�����t���� �0{��9�h^����e\��SG[;��9�2Z[��X}�"�,6���>9�Ͷ9<Ј�m��bYL���*��C+��;�>{�;�L�nikC[�+_K����M����U w��1��gQ@�`J�����:�����z�dMW��G.vq���,��COaX+�Gg���vt��b'R��rd? �ܺ�����S�w�s.�T�Ki�~�,���\g𖥲"Λ���	�'�Yֺpi����iBR˽
���
ə�c���_W�d3��&Hxy���"]�2R�@�G�4K��*���mM7����p�S���H��a�Q�����wh��kB���B;�]^E����Jc,�8Cy����PVi��F��?��O���jm˯XAd���{t}� ��E��{��m�u�/ ��K\6�uo}K��3(^m�FF��~&��@�K#g}G����F����;kQN�V�k�0F>�2����2M�x������q��g����?��R���fV<"�X`R�C�%��x�x�XQ�xN�c��hu�6�Z���}=	��6�צ��+��)��G��ɇ4(t��A�,�Q�q�8���Ԏ�6����g�7޴�NG�ƞx��������ăQ{$�L�y(�S�;Nc�r�e�+��ix��[:Ys����Q@��%�{b��DWeʴs�G����-�ϙ�͹MX)� ���x|=w��ʴ��'��;�q�B�9��v6�������I��1Z�������&��܀�Q�
��VS�H9�#�:8�*���H&ګxdRP��`�ĆJ���ܹuevE`MH^p����a�����ɇT�~J��c��6�4v��Z�"��d�n�[���E�<�3� �=7�zr��䵏IH�� K}��R����R� U!L'6i��'e�ʬ_Ub��HdbY�����[ϸ���J}_��vw4��r�@��^L��!L�]bV�y��;�[f�5�_C��OX)\�%K�Tg5��Ʃ5؀;�j�/;����Ǉ��\�5���l$��\��(�mY�}q��@���yf��k�9����Ԯ�[q�/H��g�	p�@;}o���I�'}��)1��>_�Uڄ)�$�W*�^)<�^��J�P�$d%'�������(Pȇ1��K��"�P�p�R�	P4	t��n��nT��O'f �H4��B��SF�z��G��Gm��T��Bd��pt�N'�C�8m��0� �;���zG�'��cJ��J���N'��H�`��S�\VX�o�C4�6E+��L�
?,7KdֆV�N�v^�b~	��'�iق�<�E4��~�%dVN�qx�[�b�i�[�Z�zY�n��[�X��#`��׭����-��p��O!��n/Q�_�P��u��&��(�;r�_��w�U-_V��f�n���X�^�8#���ݪ$�l�*�l�=�;S�U��C�SUWM+���)�z�L��_�cAK�ba�ڋ �^�	?��87}��h���w��f��G�"�:e{��zY=��un���kv����	�����9ˬ���؂��2����>!��A'�Ͱ���gѳ僻�Ľ��{ͤ|�[�Ξ P#M�$��{,?�af�G�F��:��+��3)p���,c�R�B��>&r\�)ׁK�J`)��7���]l��Q����h7��Ua��r�O���:-�Hn����:��e'�R�PH_: dP�QI%LU-�vTQQ���SCl�I��H
���(ۋB�;��=�2��v\:]�o�������^��Q��hX��@]/�S��ryl������8�>Q?� _��@����!c�ӳ���A	�������S�2߻��w�����>p��S���,T����p~��6y�;Tx�ԇ�[���c"��Ù[�w�PU0��N�(/½x���Hz��:io��$����&|���M`�|ec]Z�I��5�����L�ǚ�Wy`<LQ"�_8h%=ݪ��%�X�и�hsS�ƻϖd�F� 9U-�3xh�no>_�y�%� ͬ���(L�r���VH�L�����)���{5�.`�7xè��j���H��[>��~��n��u��D:��O9~ct#���yU��V;/�~�~�b����$õHi�;�&�	�H^9�n�v���Ean"�k7Dn�[�+���ơ#J?�鶥9{V t$�&�r���{�?_}��1��1�J�t?5�m�s<�ɍ� ��_�u?O��&�/�8f��9�O�P�G�|������[w-�>�M*S��D��T�7'������%'X͚��2�F/z��w~����m�|a�n���?�����>���,Dk�uJ5�qO*�gz߹�ѹ��W��#��ɇi,k�:��[D�Kj<�)OLEx�"�㤤F4��Bc��1�0[Q5��4L��e�^7���_����?mg�REbER>�w�bDz�Ė[�Wr�Z��C�$���>��J�+���٬?�oIq^��v:%�7?(#��lh���|PU�2,m�����c��T��G����Ѣ�C�akD�Y�p��ܾ��8af�hH&� �7c�u��$�޾��迗��z�j!�!��^�`����:�и�tC$�mY�d��CqT5�$�u1�_d%Y n�䝎IdN���&�ex�M߱�rk~��A�lŜ~Ts��&�GgFd=I�&E�'HBg�����(r�-�[���K̔�=���65��JR��;�k5yAϝ�=]�A$�f�X��rk�z`ͼ�R�I�ME�)~�l�<�I��d�.�LV��#3_D���Jy�&V�[�m|� �y�����C�����"F���C��;�N+u�Z��Q�H�ᄷ18
� =���hk�  �3X�^���f-LǷ��L��p�E+���H��l�p9>ǡ7|՛P�ȁ���ਢ�:���}
���o��WW4�.Jp���ߕe�i���xO�8	*�n�./k��jH�1lt�������D�CG%��Bn�C�ꅉ����/�=f:�<$]��Q�2;.�|.��] �i���z�de{A���X��4�E�}������y�T/H��p�P�I���4/��q�Iݭq�%m$T�GT��^)s��{�:����L���#Y�0��Y>�(�ON�<�ۺWU�ĥק	��90m+�]̚�}-}�=��������!����O:�V��k�鄼�&Ȍ�o!��Kl�4IF�0�,��y�+�ZȖ��Y]U�������!����o�.��g������.=��b�%-R�B����n����͡���*A �� ��@��Ѥ+\Ƕ��+q��M�RB�0Rl�W������n` ���'�?��mݪ�@�+m���i���P�bf������TQn�ͯ0��֯w����*Q�,h����_�}`|�ۼ�7�H��i�	���Q��wj��F&����g?g���2��]~�.�p����z8��y{Y�VEH���H�P�����s�Ǘ-��w�Ӭ���vV���`��d� ��.�Eby��n8jeZ�~JX�M�	��UU��QQ���N�i��C��!����*hWA����$S��ʲ���G�BJ:P#c�Xaj��[%2Ux\�Aɝ��l)8���bO�
4�� �DY/4O����=��I*���F��f�+�����Ī�#м�θ���]���*}���[+t�R^
��Q�(�a��b��o{ �璽��J�	��57��	�2݀�$M� �:��[=u%�����Ý!�����(j��9�6��X�R�/�D#CDǗOr�),Q�WnN����*|\�zK����qlڡ�Oş2d�S<]������B_��'��	�AM��?�� ,J�w�0�p�B�{3����|�jt��B-WG1�s��ys����K>!�!+ݒ�' QQ,���Z^�:�c*A5�g�����s�k;d��Þ��n�?9�����.L��2��ܱ!2�l��ǹ5�ҚX��.�S:fD���1`੮<����
EZ�_-�hF�j��Z�z���yO,�M�o�4�d@/<@��-:�磬��W�MA_�SӚ��מB��Gb��<���<���3��սj��r熫��L�d�y���ɬe2T=�W웲���ސO=F�����m�(u1?�i�U��:����	h{�YN�.R�lS�K�^��9�{[4�?�qHѦʔ��2�LYl��l2#���u��~�]��|����m;}�nyߘ��0��OQ�Gq׃{C�dmN��;HGW�]g�w������|�9��=5te��[�Ht66R�O⓶4��/��D�ۤM�����Q�5~�V��4 1�'t����57�R���_�fo*H�<��Kf2����h_ȇ�h@j��$	��j�*�r0�f��z�Ki��2��:ʍy��7��!j��nT�KpP�[��N)����tV4!�-+��l ?�e�M�Xl�;�ܣQ��K�f��#9��?��I�q���F[��7FB*���h��w�h�l|�gO5[��c9������WQ������n�?�iD!����u��'v��A�v�G܊�����S*ߎ�WիU@=�;*�)JJZ���'sς�"�z4'��G��:�^xz��7��D�n� "��t	/�!Q8SBCf���D�o�L<΁�m���=�\��.}5�\l{��n��J�Ʊ����ľ�㇍L@!V�S�:���bI���Lfx2M��)�"B�#�@i��# ���i"��PO�3 �0^0~���u���&��"����'��[���mu��?�x�u.�z�m�vE�N�K�_�<ƵL�uj+�Q~��#(��"������#?��p�8_�[^L挆�{HJ���J�p5��d�hri�{ͯ'���~�Z����S����4T�P*S�AIJ���?�;�,����4=fvԮ3�.�LS�����{�"�1Y,{�&m�M��N�j��1o~���U�Ӎw�k�Uag���l�0S ���)8�Q���o�>��!��v��UvZ��$��{�U���u{��{c�;�	�oά˫*��v�UU/�9�qP$͋HpZ*f���/��W�|�F?;��ZM��z������*]�K��Ft��5�U:'Hc{m~��O���T��e�^�}��c�2/�������֌�He�o��
k&�A�]yʔ��R4����Bd�:��Nm�U:O_ҙ`��E��7lE&�>�}�"�(�V �g璆��m����5g<�2
���>/]�B "���aE�#%xqq��>�U�t��(�92:7>�;3ه�`�)i��ﰬ'�T��^ż0쯯�Yw�d�U�r\�M����g���aqKdb{3ܪ�31��Zk���	��O�o������@Ҷ����æ��҃��T�m����#���?��c�Ne�������C9�:|09fG9�Cx��Ή�d�bL��x��ɘ��h��劒�������RN\Ö���M�5�B��ek�����f�E���h��ƻ���=T���&pQ�O���^��E`�ڒ�Dhb�6���;!�L��]㩟�;�:c�n�H�����rc-z�O����R5��X����d)�E���UY��!MT�~���~�����
�O�	62���%��T�[!���t�c�$�21�w-^nl�=�]-�y�`� 	ȩ�%��8L��s�����������q^9\�(�<l�]VH��ĝbc�7�����V�Z0ϙZf"�s����&�����������5���D"r�����@�˯�FO�Q;�%� ��|����\n�����`�{~�h�y�_	C-ĺ�D��掠�>���.�Q���3��4����!/��]N9ɡMB�]�����M��N����e���پfQty����� �]j@pk��k�ջj���%��)�m��{I�����	v��U���S%�޸��`�?��_��
�4ˉ5�	)���t.R�U��\l��zp�0��d�o7,������ ��[�u���/ ���u�-���X��o'w���^db������OЬg�G®L/�D��T��N���J�,-��4m��}�pYȭX+A�$pb��[S�t)i��]�UV�^?D�"�\��]}��*��ChV�Rh�M��eo����_��Omڐ��ꅈ�B%����:�<[oߝ�?GF(��X�U��9\���M�%.�.=$�3�����4Z�j�H^���}z��>i�����sJ7.
}\�gJTi&��V�
4�ڑ}�P��G'D�9��f���7#c����|�3a����0J�I����A����esO�"��H��g�Õ�<��OV�0>�3��5�����#țҚ}��(;�3^B[�Vsb`Io%a�Y`�.|��X�4��j,��5�h4t3<t��ݲJ�2��
._4��i6�ȴ"�?<oJ�|%��p��s�hzl8Hտ�9��o%��aRC/�'*�a��L{�I�~������8��o+����4��D��b�3��2�[����N_�̣�('����#kO��w$�Qi}���Pt�@�6
8�EN@��ۮ�2D��n�����2�EH��V�f�r��՛�D0O��1�5��0�W�1�ڌ﷨|Q��y���^����R[�L�o����t���a�=fVP}@CT��Q����}���n��h��y��$�	�b�Z�ٸ�p���k��3�j�=�%$�2�^�~�_�r��۝��8����i��A08���k'��M,c�����R�G�`�~�b����Źq��~,nO�?���)s�;Y���*�L=k�K��s0�bD:�d���g�-^|x拤?��)k�s�<3X[V�^��Z?[eչ+��fo#�pE���eb=���im�,j ����*�o��r�i���E-��>Sߘϼ��SZ�ƪd��9aVg�Mc��М�\�h��GvWg��.x���O��螚ޟFJ>r��4��o���'�۰}��r���!�͋p[�#�t��KIS+��=��8&�ٲa��ϻ)Bx��u&m�d�\�/u��=;!>��Ρ��iO�_��a	PW����9��G��/��/6���������~�9lM��B#�&o5�b�ϻ���j�,ɍ
`y�kub���f-g�x�JX��=6�7"�Ԋ�yk�/4��H�8��^t�ׂ?H�5������G��<�d���f-'������1�$7	�l��P�/ĎxܟRM���A_*�5��.'��Gջu����t���8a�	����q�C��4�x�"m�;�i���u39	�=S��2L*ʷ�E��j�WB�̱Ӌ�"�PI��o4����wG�IsqG��?Ma;����u�8~x�+�Q���*�/S�Ž���`�CcOʦ�ʍ����`Y	�Sm��ۘ�۟޺���WD:���1vJ�)�E�^ ݶ$�	w�������������j��ɟp���� �Q�v�Q�J؂8;����2#�
�s3�G"2Ű�`|x���F��kx9xe�����ޛ����#��r�{�K�Q9�}_D��Q�`Y<A��J��"�+Ê�;3���ts7�.gT�'�Ҏ�q>-����fW���䕻��ѷ����Rۅ��t����n7_r�~��>p~�>"�'^�rO��{���oB`�:*+�9v8�m�e�k0�gk�0�t
F��J�����!�v;�<ԩ��(e�؎���z5z�y��Hߤ���멩%�����	y==�N��e�a���c���31�0Ƴ]խT�A~d�f���KR\W�[�����-��lӂ��_^'aa `�-	��X�oW��ah2�R���`9������E���������We�_�O�^���M�x蝹���\SB�a��ހ���O���Gϣ�W���g	�������Y�N�W&@ϹZo'@�����s������#lr�|��fpB�� 0FZ�q�p���V��`d�'KX TI� �ztu]E�"�_D��է�|�[J#��!����<�c�f�=�W5<z}T�fK�j>��C"L�7^Ōʫ@�k�gN5����`�y�V�(�B+���
Ԍ���uT
�>�o�j��0�z`"�9>�OP��9��d��8�?&��!����(�HI�t��t���tJww��%� ݃tww73�0����~z�_��Y߷�����@g.0��z����@L^i��r1�p5�,�F�a(�[:
�E��U�´P�Ie3h����Ͷt��8yKbS34�w[7������S���R�j6�ay�^[�����ۄ�:��2J?(�$b��������t����em�й����8sm/l��Kf�l�\[�1���0x+��������.ئN�+�b����jO#"3�$���e��[}gU�4@Wi��Cx��)R#�W�
h?��I8E��xJH��Ă�X>�;������!3��?bX,w�Z�.-y���������!�[LW������i8�A�	��C���;-��B�n�#���X��&]�f��|�*G����9�Qi`!C���C��|���ROϕ�L��c_�7�?�>��}�PR�{,g���z�}^�F��X��x­�qn��^.5��)��ӽ�Ī
��$��eI4.�[E��a�	�rA���
{�D6��E�p���������.�iH������ޗ{ |��s�C�b��P�v�9 M錅w�3��;�x�T�ti�r�\tj�*����j	�����h/(G�D,�Gi����R�v`�XrZ�Z��˚˃�z�\�{-��-v����$����>�֞/a���C�M��/���ærl�8n�}�08oM^b�ꝥ�ּ'�#���d�R�'���}%���؏%`To��LƋ/�w�Q��&��4󶣯v��0����ks��Y�o�&��*~��,h���� ����$��lg�*�)�{RD��mU�S���r�ޛ,a�R����??�w�Z��)�GPy���$��-3��lV���X���w?�%M�bi�7�Sl|/�-��X�����	��K�2�B�,�꺆���vzl�p)`	mD�r��nG�L,r�?��g�y�Q_��N���R\w�EVP@�Wm��"� ��Xߦ�)��Qg��/�o.*|�z����6��g�'^�\��_��8G��\n���O	A��Y�E�ȯb���l0��R޻��R*4��22|t�s��Aq{�&1/L$r�:i��g����L��]�j�cYjU1�A�0��7L�(���!K�s�l&��f�sY�t(\'g�M�B4�_�"�6]Up7»��&��\�s��e�lK3����S�N*�R)m��Q����ǧ���B߫�ʵH5��������ܾK=DJ
�O��`b��͌:}Q<��zm ������ߴ���`z����ۏ���8�:y�'�H���N5��G�'{9�Tg@亀��3��R�����hD�37/]��N��MM�/����S�.��*��X/t�#~ɣ���3����y����0oEO�[fx=�C	�ޓ/����"g9��M)���7)G��*���>,���"`8������<ym��I�������e=�����eF0v�ҙѻ��wt�Z]�Q��=$#v��s����`\�r��ۿ"LOz��s;;�ޭ٬_.�� �HW�E4�zE k��m1��4��!8U���7����J�����Ao煗;
�nv'�<�tJՕ�$�0C�ԃ�;��^y��w��Xi[�2]�!ю�/ƭɍ7�C��x����̸��B)0����z%}h�:T!z�m�L�ƒ��g�/�����u� %_��0�K���[Gыw�4:���0WN����G����h�j��k:��7Mn������ee=���ֵ򪭟��v:]�{P�P�Y�gi(�w���v-Ckr�3h�{���}��^w�n�9�����SRTY/��/rCq�J�mE��Q"?;Q<L�d���$��GzUۛq�r�Jۤw,��K{ד3sF�G!��x�E��øuu�B����gvo�u�f�"���Ӳ
п�>{vETt��*"%�դ�;��0��M���t�a�D�<�_�Sr��zGoڃ��ЋF9���Ani�����q5�,qQ��m���igV�h׭��[�/6O߇��.G-� �=�8c�;i�U"B{���R�1mq�r1wнIp<��8��z��̇MhD�$�E{��M�T=�$n�r�K}����mI2u�DM��;��n�����ĉ��1�BY0�\{Ǉ�:���^7'���hG۷��3��~۰�X����M�(���<_�d�ό��V�ilK�W��	�a�z�<ob;�_䂟P#H�s�`��m��j�u�v]�K:R�qj�E}�.�D��U>b�QG�&�xI��4�c���Z���|!�Ȭm�ٳ��$�lA3.�̎��ig]�3kGܾ2F`vO�Bi�Ϸ�K�H�墡e���i��I<���'^���O�.sr�sJ�"�#s;��g�%3��g���5~�8x�@7ý���3�Ł��=mi�T���i��7����V��OT�A�fږ�L�������K�D��䎩�e�$��Gp�AtcT}�(���c�Ÿ���җ�ѯ��ufSh�&=�Y�aOx.q:ɘ�.�m�˿��v]("�Hs�Kh��&���q��[��ۇm|h�t[�pn9j/V8�7U7�>~螵8����������I�y���WX�L����7�3�k��g��B�>_��)��YU���W���W.�y��4낼.��l����
�����vQH����<,ꌿˉ����Y�y������"��w�e��ٶ�x<����F�_M �јh�g����xKN����^J�ӥ��u"=�\�[ �8B�þU�[+|������x����:�b!����d�Lo)r���N��*	�km��B�G,��sU$�쒐~��]IB��[72}�E��Hp�}��+�c`agpv��H姭�0�a���Q��������-��ӧ�Z��%�M~�.���������؄W�.���m_;+�/keWV�Z1_��y}c������	�c߳=�Pv����-���l/Hβn�o9)<yRB��M̧?�@,��������x���R�4���==�4�=���ys,�����Ĭ���1�A���k,��wr�(G4͟jjۛ�J.>��jX�On��o 	ew)�2�l�����(] H*H1tk�}�*����.�2Z6�ğ74� f���������ط�w���3Uo�!lS�8r��	�T5��w������w��lI����k)Q����KB�3�0����U�º`��q�z>E�夷o=��@���F�9k�Ϣ��]X65���J�~�$�-�3~n4����b����XY>���֩�O��@����d�6=s�;Y�8ߓ�q��|%�	��H~��C#WȮ"'̆ZY��1�x}��,�I�=b�P��^Y��$z�O
��ү1냪�et�����fD��������P5����<�S�~���V����0�}N�S���~�$�_UQ�P�MXl�0��&?/D��7���'�E��L��jyQw�~��]�޳�&<8����r�fG�<�P�9ц9�GgOj�}&����L�8����V�%�Dg�%��/��̹!7��H	��+W'j�9��吠�RO�省/�o/C��_��9����v���9:���\��[��l�nx���f�Km�Ұ��θ�J�윽�Zps6���~�0�z/.mX���B-��P��K8��w�����J����{�@"�e��k�D���'±��۵�V�<c?�W���t����-?��|a/'f0�)��>�F3SxAf'����4zzC#�U~�r���������&��[��d��\bnU��:�N�0y�Z'ᘓ�?�M��|�|�a��È7ݧɞi*:����>odE0������y:�~��L=a��<�a��4 eC(;:O�k-
�_��L?�Z��[X���W���j1��ʝ�|�]͡Q��h�
�߂p���` ������/�J��!��C��u�������9&����kJ�>�s��X��:��+��T�-�3W�&�0���7ǥ�K-`��7���R�y�����|j����f�V݁��'���;]��͐����
w�� �#��������GWh�m"�u$xŜ �<(��>ҎGM���\����]#*�vQ>���J%ƌ�r�Q��d�^	U��� ����H�un�{�^�$��yE���gE�o�m�7A~^˶ߵ"�;����ON���%M��_��\=T	=�R(�i��x�����N���f���,����IX}�@�s���y�"�͑��X���vS�h�q�}}�ɼi2�}$�#��y7� �}8���������6��5�o6����+b�RF%�7�GE�uَ̅�?b=�:8Ē4B)`�[`�z�������-�3[(�*V��z���b�������ͦr#�!<�����L�<�`�K_���f�V7̙۬Gg��/s�o2��TȲ��-P���_�&^u����=��P�!��Q��D���Ʃ��K�N7��0N`���k���E���숉����Pr���w����.5����Ұ2�:�#��ʳ_d0�1-�����ph�S,^�ԉ�s�M���"R]B���3t�e��<��V�Z��U���R�cmj�Y=~<5b��B�xl81�N	��G	8d[>}N�ݮ;���6f?ա\.e�~��&N6�&v���54��%�j���,{_ɿE8�b_q>�pb�8Bh�k�j������u��F�d����P��������/K嚱aJq��3]�m��݆�=�bu�6oyn~I�Yt�J1g��pr#͏�)]b�3w��Q��X����0C,�^H3�gN.��ؓ�6s@��J�h�<��OO�=
��)�v��B֏���ּ������X��-��z��}͓p\(�g]E�;��$��L�u�|3��P��穲�SR���i��C�K $�׼�3��h���u$�E�s1�{�����q��0�dF�Z���1��Ѝ��5�Cǻᦒ�ض��ű�/�-!^���M�S4Ţ	I�H|�ƛ5{O��C5W��yg6R!M���]k�%B�N����)z/{����C�w��)�*m�Yc��w�g��hv�io�����A��g1�����$�o��
�5��=��-��Z��!�|���7}������-µ��M,����lG�n2�r�.����S)GxW����g8�B�Au�:w&N*C�=j�3�Ju�;�uZTx���4��%���t�M��4}��xÞ�ܷ�( ��M �����%�ݖ�~Y���|�+�)�ꓫ7�Q��G�a�Iy��5�����5���}+eR�x3��Y>R�D�p?�M-�^��YNUO���z6�%+��''#6�[�WW>�4�4Y�,Y�e�)sYC��3�ظ�K��i��X/�Ev�f��c@�P�������O�{Ϸ���'�Y�4����qsd~N6Oܘ�|ˣ]@�{U���\����e�]*��745�?���K��n�.�ѡ�|"��������rH�I
��?�z���	��O�Tv��Kx��hO���0���nI�,�Sj~���m��bd�'{�sx��i����5���0�9e�3d��L�%,�>ug�Ӥ��β	�<��@h����^���$<d�{!H﫭Vq�����ل��Ek���}N�"/#����{�Λ��P�7�F�X��_��&�QV2�������'�z�܃x/=�{�#�7d��x�gaΉ��7+j�C4љ��|��~[�u�a����F	#9~�4���ul�{Yguf���#l3q�X�x����K؋�5��id����#/u�H(⟯�V��7RW�$q>m��
|��`�E�c5�W����ջ�6�}��`�����z�W�=>k�1���p.H�R��y>3�IO�VՋ#!�s0=ش�j�}Ӻϖ���r[��&�z���[�Z�+���k���v2��왳o�l�� \Wi{��i�y��D\7�:G���'��d�:Ud�|"�	���SQ�ýoӬطx5�%aZ�M��q�I*c�?��!�e}ڹnHӱ��n�פ Hp�N����v;Z�]+2����Q�Z� Ȟ*�x)��`λ���)j,�q�hj���Id%q�-���_5��\�'���^�(Sԕ�?��^Z�m�Zq��_A=8Z3�J�����kH���[ʥ�~�yF�j�o	"���N1����r}F��;��-S�Q��d^>yu3�	io��[x���9h��������r1�s�z��eMOO���Y�VI�aj�b�!�6�jkJ��@��'0y��H��3zZz�|2pM������$}�k��~OPh�u9K��J!���˘�ߦ�B?~\�b l�YEJ�N���|xo�W����"\����82U�[�[*2�Q�΃^�F5A�Y�U䠵�"��~_g���������S����Kt^�ٗ�N��d�w�#?+����@}�����8:4�h�ѕ �������o"H�$�h����.,��5;���,֒�q#�����>��E�멑}�$��������gg�_���ࢄo9��ަIsp�\��]�[��UT�qx�KAb*
�8>F| ���:�4�l�J�}Y�TgB|��8j�����Zu~�r:��s-0۾\K��������ۜ�㫫m.N�C�!�Z$�����~�}*�{j�෍��|ͳ��V��9;l� *GMW�y��=H"_UC50�tl%nK���{0{�^��sOƼʥet�nɕLr4p�?�: �c5��+�Aۜ d��*˓vh��VNI.n`�jae�����5�Xc��.�nO�c�">D�G=���e�\�i�>����������a�\�g��Gk��Ⱄ�}EA*��p[Q�=]u#�.j˧+���5�2�\�@F�F��՜M{���v��"_;�K���$���n�N ˎUQ��!�l����Se�����D�����P� �!����ye/n��S诣��7cK�a���#c�- I�_��{�ر�cnf���VCI�]��F����K������tB�;��[�/=�H��VW.��ܫR_�yxu� �V[�]X���5��_�>��'�MU�??G�nd�-����~�8d{R�_�����S1���:cph	�W�G2���Ԭ��A��g;Tѫz|��l����Ys�I�O��|������?"+�j�}����-\�5����{�����s�n���A�%��VT���-J;��F�A|;Q�,x�X��|7%�8h����^[G�LZΞ�p�EZ��Ȉ�<�H &)9z/�{����f� �#+�'%ʃ}l3����}�JK ������(-�tOi}哏�Q��+�ő9�@>ވ)Uś9�ĿW���`�����<� `�Xgi��x��?Wn6�X��3&�}zN�+xr	��^�׵(�sσ{\t鉳ʞV��hkz;�)��d�.-&��:�N|�*�>�K�=B2��lj���N�uTֶ֙@�+���|﷢�c�O&����Ȼt�F㑑����SZ��/tVY�~8_�BSj��Ν�5�w�L��J�G�;�u۴<��3���:ϳ��֮x�z����>�OzQ��=U�����1�����F[�N���{�?	�|ׅ�J�"��(cϚ�I�&?���xᡠ[ue�x��������$��:���C���b+s`��R8T��u���"�*��n��@�T�ˀ�+mgֶ?�xp̥�j"3Ŗ��+��w�b�ˍ>�Kce�V��,&�f���C�l)lx�V٫���l'!7B�����5��	Y�F��"b��K}/"&0�|b�`:�KVj��"(��J�]��k[��D(�R�$���'����I+�P��߳��Y���`�M�P/�l��H�2����y��)�����Kz���B��:�6�L mݵ6��2m~}��oJ��0y޿�+����r4!M,�`�u�q�XB�V.��u�e�u�l>+��z~�\B�����qMc�3{���h��E�����
��p���'f9�ʅw���q�A4���-x��^n;�,�y{��@aQ�#�h[�%�O�pn�iP�T�և����x�����sF�������'�W]݊�^�z]�J	b�&xE� Ѧgʳ��[�8���5��4Z��$�G��ק�99����Z7����}@ΐ�)%"�Sa�+��>��N��0�d���0�(���s��CϬ4��e�B�����4�+�$M'u9�x%~�R�i>�=�U~,��鋐��Yn������,CN�����{I�rX
�y�&^�X���~Bo����FPl�D)������}cm�sS���t|GS�����p��M};&�����R��s����I�#��)���qn���s� .쉤�v��4$^T�����+�Z�^z�0 w�j:5�gk�sd��<��{�!l�(E�m�p�Hv����Y_�l����Snjog^�^<�z�c���%��D�\f~��"�@�ֆZ���P(�_a!����9�U9'��&��${FFU 8��\7]ז�p�t¡*=���1Zg��ko��jK�s�\�u�Poz!ۢ�ǍO�c_�z�5���n�	z�*~���,G�֎H}�>ť�3b|��{'�M/�xo`������f9xRe��N�����qt�+�b�*7*�2�$}�T$�b�k�	 ��=�YE���e���[Y�e���+}3�=��'�8�ٌ�ѧ��E��>�9������X{[�d�5����z���U���'���T'魟W�4l�ږ�dZ,�\	X*I��Aj�����3�G*ޟ�NXXT�_��*&
���X�ca�P/��(�}m��ڥKS�5�>�jY�م�f%bo���ܽQ����+ 7��i�hM?x�V$�`r��Cq|�p���h���Q�m*�����]A8�����Q�dz,p�n��k���@�#ă6}�_i����ZXKGxgF$'�mɠ(Ϸ�Z�2��A�f���]�{!u*"͙�`
�*��G+�������ic���WW"�G�o�L�L�|؆��M924��TKY���3�����(���+�a�\S�r��Xhi� }���a����<��*������;�Ǯ�b����?<E���f���z:7њ�߿e�ƍ�<@��O47�r�A	�"�>ș�`�����Q%Q�u��֍'Pj0-�4�]�m�iC�����r���'�J�!m�,ȁ=1trM�ʯ��K���xop�TR�x.#�m�Z͘	���vn��gY�}����zw���} ��z�\i�f�QU����0�b�\��w�5�1�����O�]��0�kA<s�&i��щ+��P>��#�s��#�m�Pdr�;�.�-��5k_>K=ܩ��f�p�ds�z���A<!5��_�?E�(�,�4_�:)���LE��8�6^v�P�Hh���H-KR'q��%����ha�&�pOj����rf˱Y�hr6�줿�7��}��R���J!6Ŋ_�_�?�qGO�S����� ]'z��X-��	�Y�<ċ�#��p\�a�o6���)�m��e��K�Z3{"�}RB����Đ3
�seH�fe��gY��կ�E������5��0=�bX��I��@/�����,��!�����C�5Z+6�4}8�� 	�{�������N��䁑&�z�I�"�K5#�eS*1��d7��z�2.��8���\��/Hb��3h��f�"��d��{�Q��=�ũy��&T�vx3Ǒ�]_�`�����;h �g_
�
I���cU��rª�oZ_��0��yŢu�&vm�k ��n�]q ���a@?Q.\s���Y�W�+���+��{_�w��:&��x�-:nEs�"����f!OI�����ʆ�S���zRd��R�������+�Ʃ��Ɔ��׼�[/7�rg}�'�(�f�n����(C�4�,��Ϣ=1߆�V�Vt�-�΂�u�Qi��V�T(��w*��ͯ���@K�����Bx��sv�t'����aN�ݤG3f=��bv^�!>}��[*����o3��Yd�(�K��WS�睷'��`����
!��r/N^��s�DU��!� �1�����u�sJ}�����'_o2*r�ͺS,\
�j��f%wGQ���3�'(F8Xd����&M��M�AK��}(�ᛩ����]��z�ɺ$s~�k_H+���ly'�#3\�r�*y�.�:�T�ԕf��+T�㉅�瑘��h��c�m�24s\4�<~s�5F��T��S��`Jl%�2ZI���gR��x�����x����Nmu=3����0���~<�X#���,ph��XX5�T%�m��f!̚����C�}f������
����~qOe��zdݒW?�|�N���s��;SUe�r���D�ٛ)���;Ko)�h9�e�DD��0��lޖ����2�mQ��1~�'�s��[}�Ň�����pm��>��+sWCp�w�'b)�#TQ%��w���DM~⯂r�8�X���6���ơ��D�J��w�>�H��� wI�����ϟ����R���Y�ܮ=��L>p���:���xGWdudT�dl�E����u�itHBb�qX?��<�GRs��Sv��	����9�Yx7F{�G�F�9X��3=rH�zk$���;�����\X ��k�jܴB�f��ɶ�X|�#�w��p�'�p�y�G�.�GC�9X�u3��_Ge��Wk	�lֳ"�=T���c�2�)s#[�ݎ,�z�ξH��e�V�4�2��#�"��$���_�Ԙ�@��U�!�j�8I�p;хi��7v`����&����n�-��[���7g'$6���!o�Z�D�M?�$�y�<}ivI�+:#�[kklÄ#v�g���[M�1?����s�y�{�����hWt
�
��Y<�v7�r�������.���-	�,Gmnjs����|�6`>DHUhJ�5��&@����[T��0�8(�W�Y7����g	�IR!Hv�.m��]�;s)�W�6�.��g�\[dD�D,w���b�N!�,oPe�V�j�'�\m�;�l^�=��������^�޸t��!��Ɠi�~�g]�M*$�x3��Ñ1X~A�LPF�kO^^~|5CO�B�AFv��G첦qTL��
�>���:��U;�T�e��
 ���'�DA�s�7媪�.<��	]�4\N��m쭒��82
ګ^OW����S
��,0%M~HHd��x��[K�,����S�1�Vy�̌��-����Uw��E`S��|m��U��S�J�Tn�d��7>b�Ga1���5��/��Zt�û���m��]�M\$�Z٨o�<�LK�;������T�cR�嘊�z�����]�L(��!UW�l���(-��?`��4�=ۜ|yuumQB^pi �v
��j�Δ�\Ս�3)\>4��^��������v�����,������t��hQ��N(�OG�#e3�r���z"�D��� ��J�q�n����h�x� �pl�z���i5�vZ�qt?uHEO��U�].�-�LZ�U�숄%/�K���D�]�����JmN���I�:��E���6��,��/�w���M3 �F|�ytT氄~IV*hX�\HJ��u�N�̃i���}�]��T����y�Z��?����9w�D���Ќ���w̌�@'/O��\�7e��ŀ��V�$S.JU4W��S  ���'/���Q(���)#�j��3d#l��%��1�tu9�j5X��ȍV�o��8��y�.��A47Hh��J&#�"Q9�!^Yf��MV�$��oj	�]�3|��>���C�0����Y�.�D8p�n���}���Nq���;?~0�!�H��2�[���ǧ��\`Sr��U�������̏q����zerR�.-+�8sZ�2^�i�����X )~��>n�<���]�=[O�
1?�H�ԍW���L��,DM5M�ǒ�.%���]�%�:�o�_|��۱�ɚ[^nk�W�U~	�G$��^�2���q���(�5Dg��t	s��l��ӎ�&s��1�?����965κw���̨��yY�e)$�=t���_z�
��P&\9J$X)W �K�]Dƅ���`��)���������|�a��=�;�kRwiKi"�om���$F�&z�ݩ�Nic ��Z����'�E
E)l�S��Pr�e�Q����?#�S����2�~�o�9"�G;u��Z�/h��azB%aEe?V�k�m�I�̳ȁ9ú9U�E�K�a�rh?�b Y��F/>����U}����]dH�=ҮU����&��7���	O�6\� 4����^w�1���J-x�fp�4����/3�(2j�o�݊C���4DFh�� TI+����K�]9J*Y�3�qw9���ƫ�2M�B���o5Zu��8�Ց���<7U�Qo�h�Ñ��d[@�r�*�[R�5��*���ȼ�O������E[�r���`!�䋫Cv92�]�YK7a�:��
����~�������{�BJ ŰU0DB�]���t��h��b�����+փ��!�?�?�bR����u,���K�v����0��#˲8J����V��e���@>�����F�^�|����:F�r���~�S������͌㨇�ڧl���V
�mV{H���M�5�,�tpq�:�74�t�s>�|�b�P�Jk��y]/&�?�������9h�J���O����������W?���n�/�~�ܘ��T9�厊w&3�=�n�(;/+k�V��(�<��.G��]%.>Ĕ�
;Sp�mw�/���sV�r�ӗ�(��tM�'��Ya�9�b�#!!�]�o��Wc>���,3�YOJí�����*X��Φ|���sm��͈�}���ы髄��/�
Ķ�b��"�m�������
���n���oӡ�y�=-��F�"�g�����/d���%6�����(�z���hU�Yr���K�\�,]v5I�܅%/�+�~���0Լ�8L�|���}�E���F}C���s������y�-֗���9�$��<͂5�<�/X���+-��t��߱u[��z�ͅ����_6f�����w�5>�m��r�����X^��i7˥qc��r3���81l{w�.B������w����8B���/�qց��\k�d�'�k2����*--��^���bv�Ȗ�KM�F���������p�}PU��m�Zcl8�Ѐ��Hl�d2~e�"��$z���[�J��/��buL�{{�p%Y%(0�O��5-��}�?$����8��u�<M
��_$��T=u�×}�I�@pNؔ�_N�#b[�d�i��3q���4�O�=1�+�f�#��N���x ����~�I����ܟώQ�E�4��u�����?���<j�䘧B�2�!BB\Ы����9�-$�6z"�f1�����g�,�ym�'�t�bVC$M�=��
J5|��5��K8��X8�wm���7���1=�<kv����9G4� 1�W��м�f��ȳx��9P��^�^Q�"qk;�\�{���)�r��E�eԌ�]޸��3#���S.ӱ�(U{��S��-4��)�C|]
k&|S���ˍ}��lo�h�$�^�Nm삘GXx(�E-���.�Г?S�,7Qn+�A��r����ȴ43�#g���a�(%��!SO}�����x+}��xx��&AC���l�PPe��}h(�y��UX����F9+$��a�h���U��`����
7��NT@��)��r����Xж��'���'k�s.�)7��^-����������3�+{���dB�����Q����"���H�h��8m�{����\������ɕ�+mc1��;��mng%�g2�}:��8�'L�[��Sa��B���R'�W*Ů�J���|o�4�PX'�����.|k*,)Qӯ	���)�15���I�jdr&ڌiW�6:u��%.,ݭN�W曨获y��f���ĕ+9R���[���q�C�4�
�'�+�(�7hƆx�n�:'�$����׌�F�m"4��C��;�{�Y�n���-���ϋg�Kn���۪X�fQ��԰������f���f�ӷ�)���{*u��鲰.�h��kk|�5���"]�F�Y�^�y>�-˥mzM�F��� ��_�g{�1�&'1��旾sA��7�N�"ɀ�o��iz/L\���M�y�Go.u��ʻ#%�G���Z��z�*}�vp��&~xe�.�b~��;m�M�C3�x�C-�Pu۝�W�"��'\S\�z��&F/�nՓ�x�TYN�jG64롦s/Bf��iB�����q��Ƕ�� `���Y�x��z�2#�{<��qNzt�2��c�`T��s���g�>m½B�Mf�+�꣊O�h��.۝��v��!I�%־&��7��e,�\���V�������p?�N[��$��\�"���v��h4�~�`�q��=����N�P�Y��/!�v�5٣���z�ez}��M�(��-^��my�]�wc��[!ޚ$�{S��<�o���/	��/���3���1 ��C��[�a$G�#��knw�r&�7��)j*�q������Ť�� '�����}55Cf5̳/7bZ�9��Ě��U/J9 ;��B� ���� ��Cz˳�_��5�N����+)[dYC7-�nnc�:wv�;Dnb�k:i#ШM�Yl��| 3��4/)V��)�5!��|�KV
�Ȳ����������pR��r"����Z��C!�΄�(З�͢���7?��F���z���Ug(71ǜ�&�r0b��i��:rYGC�W�ɻ��O<��?�[[ !��j��D�y"�BS���+]���ZE/�L�DK������|]���O^LO�t�'�q�^�l&S�-��sV�X)X�f���pu���k&U����=�o׃>*"���/W�c��8֖����"��� 1vl��z.w���W��G���pF�T;�t�\+�H*u�������[���l�3rP5 89���bm��� Xp�[���Y;�gKlr��M�r	��d��W]���3ͧ�����[Y�mn^�Uί��`�+/n!~d�'X(�O1�Su����T`fP��x�<�4N����mA/VW�h�x�&�Bb��3�~�N6�jB��ƌno��6[��E��\�!���/ɝe_���h,�ƈI��x��i�߈�b�mHh��DYPP��K������sK��чľ�P������A�P҅��rV!��K�ioNG=5�gs�Qhh���'㬒�ͳb���m_�(����J��i�%*͔F�f	i����"wr����Y���ڎ��ԡL��m���e|hH�񶶾���[�b���0��Uv/�d��ΗW� �����+:��n���=��};�N��YG˧D�����S�b�Uϳ����'��B+�����7��{p�,:W0��7�������9��T��6�y�2ֵ�b4g��G| EG�M\�\G�������/�!U�h&�cMy����#S���;�|Q�҈�iv���&�&_K��{'��d$�}:��}Ǡ_N��8��GS6�c��ʑ4�%�EӠ(iM|��kX}��yM�r�4�qVF����[�Az�}'jy
��4%C��AY�,��O�o����O�v˧+�z�	�J�����u8
Aed���a���1 �+��᥇��M�ށ�c��/��R�m��!-��b��uN�lc;k�7#����8i�e�m�JA�����h\�oӴڦ�P���-?K	5I�d�f���@���-���@�t�qnw�G%�|գד������-ݧ�����
�%0]�+[%1�����εv��n|�ގ��U�^�U �	B;3eR7:*?g>�}�u�<��˺�����	ā_�J�U����k�$�4l��6ն6gԴ���1+�y������ǂ�=y��k�\G �pǆ�f�˼ſZ����n�g��x#ȟcW��x���p�p��ɇz\r�N��K�;�F�y| y���4����TVH�TW�8�؂�,��f�ț�>X�,���������r"��[�S��	���%.m���%/ϧ��K�pj&�#_Xu��u�â�"�R�}-�Y QX(Mݿ�تm�����`CQç����p�"s�9<������Ib�jޓ^��IsIڬ�,J���6�K���M5�c�ω���3�_"���d`s��&��/�ʟx��E'��<�5WZ�s|�>a�ʮt���]���k�,����I+���VP�4B:����1R���XJ��r�.,�b�x�
�5�˖��6ꂌ��.�G��q�<�?5�H�Ev8`d�+-�B�<��H��8`v��|e*�s,Q�p��1�3=��!���}vz(.���`���$;�Lx�hL	I~MbH[����+��^߰==%)(J
H�Q	i�fJ���c����ь��3`�FH��QcCb0���>�{�����~�羯�z���VW7�:rU�+x��:��b�b�Ɖ��5{!vP�'K��Q>.�e����%�Ek�S�A�ÊW%�_�CLT
t�_��E턡M�o����	��F���Uw_�&�|m����6����4��ܠ�us���v��5P8��{X��?L ��&0�uxԚO�U�C�nY�Q~X�����~[�V����/��;o����=wpT� :k;7���6} A� �*4��[����D9)(��La����7i�B�n@q����\��0>�"���Q�j��Tg�_q,���;ͪ)F�r�Eٌ�>��p����m�E�P�kT�E;�v���6tY%�N��N��GǮ����ue�,OZT�%U��x���=!ϧ�x'2���^�?>Q������	�b�(j:J��a���@zلW1�U�SX����N������]��i׽�Zvz.$��rJ�e�i�� �l*�1޻=I�R?Ϋ'ζ���R� EQ�Y���� Y}PS��bd�NNN-zq����-)q?�r�G�?��\A ���!O����)&z�].�z�_?�H�%
*�=r��>�"U��}���u7"ɗ��� ���na=E8����<I3��ǲ"j��0z���N�q�?���-|��/��(UuO�I� ә����C��`��P��$G�ʕ�~^L���?�_��Ljd���S���aa�C}��ʠ f����vv������	�=�?�S��d���,C��O�� ��xaX^zV�R>"��7���efT	��RL����o��?��}��o
Z��u<������L��6�Q������o+2�Sf�cSW��ӎ6�3Sk+�>��a�[�2�͔��v�y�S�!�����c	���p�����`�WCeq[������a^ �j��8Y�9"��#��s�=�(m�C�*��;/V���1�>Y��it����RN+�E溻2a��h�S�5���׳w�D���gZn���ތ���L�i%������'ps�{1�<�� �ء�il�B�8�"ۃ�z�������c��ΐ�Q��|MB&�u�}����r�dm���v="�U]���,C�g�R�����qs�G?�ɒ*�^P'�x	t'S������'д;|��{U��?��z����F����{���$��I��V�Y+�Q�:�������O)%�\�n��[�.�@�v����i���8ό���ƾ	�{���騵u�C1hO�ԋ��c�(����TFZBC�5�'zϭ(�[A�xP����|?�Q ��畟�sr���_�y?#g˗F��L\���V"����y���[z�E��=-��d�!�e����� ��PLo"3�e��>/zǀ�Á-ŗ=V���6�Y�#�נ���!��m�S�S���9@�Am�Y������|W�C�yײ�.������|
�YNx ��s���l1���J����J�Z,n��U
�gG�t��f�O-촕��J�I%g�����
����d�1gnJ�g��ۉR�F�9>�E�����U_NY��%k�2�:�%}�H��43�Q� �}���s��i`�c�W�dP!�-s%�sP�}vbK�ה�(��� R33�a�k��pHz������G�O��M8�-Kɞ:����pD�oK�]->�,��� ¾@�5��y(���/1�����.���K�d�Tغ�6�>`�
�sy����cC�����#|%t_���I��Q���ƾܘ0�W��M�
<G�w]����
�_����i�Hx��G���hQD�62*�ef�\k��{ވ��q %�R;ٛ���H�Nv��1��KQ�� v
W��_Y��;#���+G��+��9M�Y'8�x0�H�@B�[��+舃;c��l�[��(x��޻��NѨ��޷2c�����[���g����H~�rhu���w> ���rM��O�����g[����@�z�x�A{���N���kC�FS2(�0FD����ߚ�ۅm9b��+�����RyQݓ	���ó/�*9�ꐌY;W�`�������ڪ�J�$�Ҏ��pt�2hJgWQNP�"�n3}��?[����=z�����M��%ԁ�x�ֻ��r�����!G�����5��E~�^B�8_���0'������ྪ��>�������I6����Ш��0�������Q	&�?��'bCF�a.I�.����"����>��|>�6�2�{�����4���X�M�*JȂ��0��U���^S��VU�2Oe�cA�u_��i
q;r�����3%��<U\��ܼD�R9?p���2��'��\�����W��4��%b�zG�B�a��Fpgnj�����[�JF~�����H�U[]��������t�	�c��[���G�!��`c��t�pi�Olu.�	�|#��%����P����pL=k�T=��$�(茴=)D��\��;
��S��z��z���3%"��9��,似]-��.��ZP]�}IT�ճ�#��4�/�q��k9s���#�9�B��A]������Y��B��GJ��Y��)�๎�c�smbn�Kx����,j�0(b>�ڼ�x��z-mՠ�_&������n��;����M�DQj�g�5��$��h~5�����U���w�YZ�?��1,;��u�Ik6{��5~�Q����+%�eW�:�y'�6��v3�`O�V�6oz��@W���?������p�ކ�T��1�I}�c�_9�Vg,�=V���K�L��oA��lk{�c��F��e����L���q�Q������;�'$��7 _d��T~�@8>p��\��R��ދ�	YvM��Ə��C���&	�@|v�s7z	rneB��9J��#��>`�z��w㴐tg��c�Vu���$�[t��Ϝz���f��MW9�:�	�R4�涱�Э�"̲چ	w��Ӱ]��y����)��^��zX�(Fg�`7�EN�����әl�)�4qL����k�J�s�I��,oQKM����/��f�y��:h�~�y"��l����쟩�v�Q���%��{c]7�o9We��Gu�	�������#�'�+��O7��$
����T����m��6P�Sn)�e�t\Y���a�R��<�O�}f����u1w�}1��J�%�'ٵP��AqԘ�����A�z���`)`R��$�j=eS�ytm��t��7\#�g����y�YfӬ2���9h�5���I�gU0c��tvb��)���$�T|����wu�ؓ��;��L&�%��乃̢i!�R��!��?�)F��8�6j^���M�Telp����ie"����\�c�y��q����D+P��7�����/Wp������ͣ8	I�=�� ����ke�*�~?������	��쳺:��o�����7H�RJ�)� ���/���8�Ɖ��kg�[$Zl��LI�ȧ�>D �d%ʗ��6��:~ N�=�'�o�<X�R;�N��;־�'-�b�A������O����4)��Y��E�w;w�u������߇��q�N��x2>������(�򟆶O7$<�it+�N��1~���I��2��2o�X����[�%� `�a����(�-1D�W�;�Kɴ/����ƯY���������J�@��2��$�ï�G*�(q��=��ٯ��g��?�׳iK�:'��`L�3d�Gn��v�6e����rmh�� -��i|9嶼͜�Ω�qu�F̺$ꮖ�"o����������hZw��tlV�D���{Ͽ�?��ͻNZR���_��!cq�5B�G�-2'�y: /��r묹���w�>C�W����LW����ˢ_	�e3\*n�����g?
im�/2A©g^����8N��iK�ծ�_��ćU�H 6d��#ݞ�T3NZ�b�C�_c$�X����toMRC�Q��{�����&h�Y~F9m�jw�]���Ͳ_�'_%bR��l:�Ӥ�M�8�.��N��ꮯ>i3up�C�����lӳ��J�}J%�9$c������?�@�Xk�㶓B3\�S<�OU���t
��������4�4l��w��I��X��Ĝ��6�-C<p<�8C��0��C�����P���y������&��#�j���jԼ�����:�QĆ�x�jn����^�]�� }�f���y�(v�N�D�K7t�~GO�����o��ԯ'�WO��e�,+}�53����nc��w�G�.Y8��yk������3���>3���Be����ظ���8A����R�?rH�za�E1����#g!�H#��q��|�D̫۠2�͵�C��oj��S�Y�,Թ��@8�nŜOS9�M!QWJ��(O��i(��7��;�_t�*1��S	�o���\j_���R�3Q`g��VT}�ў=��fޅ��Yp��:ب�7K&�B��!�h��ʯ�)[Q��C�i<��W��_)	1��ߝ�K��|܆��m���H���,��Gk�J�瞢��<Q�{	�L{M�>}VB}C38	��F��]q6'�El�En�3��?�S�a��=!�?%��_��4В�l��ض���Q y͡jK�h��n  Zcq6li۾Pk�K���^>��ᙧ��1kq�;�Z���8��aSwIc��OZ��N�ކg�W4���|������Ž�?@e�VL��'#�1����/��dU���g�)q�-jCOl�Q�nh;Uo�q�F��T"����s��n
����ٴ�晬Fj�$ݎ.P����"g7����6�+^̨2{<����s��I :��f�$A�d�*\>�/�[�T�d���4�^�'��v�����r�_�d�V�R�T!�]��{wO����4����?���-�L*$i�f��4�N�>A�j�*U#�Ȍ�D�@
2]�tv��e�\�ũ��亘P�EJQn��/ճ�K����)2���J�pA�έb��vZ�ɱO�`���fJa�=H��4�/��ָ�7V^4��P�]G�&�M�
U%����#��G����=N\#����N��*`�Č��_$��1Z�@V�R��;!���@lAQ�R�ٵ�tW����z�M�P����C��W�}�eK	�8ɫxW�@`E���2p�4��m�6T�j�f�%���X���䬲2��FɁK�/�G��̖L������?8���[ӰY���hwƺT��Rń��R�[˼z��C��?^�^�R�P��j�O�	����x���*y�,Sz�l�KW����j��"��yE��������rP�kD����Y���z���k��:/!�"�U�Ze�[�w=������:M��Lfm2���`:�3� i�q4ӎ�¹���a�>B��B��g< �(�y5��E��$M�o����/A_�����Ļ�$6��J�����z%^��v����e���\&��Jތ܃3������l�Yy?:}յ��08�w�U�݋�ɫ��f�o�o���w�5]��,�_M�D���5�:7�r�"������4��}��.);&�V���x��"����㴑�| !C�_�>�ո�����?�/��`��~��j�"���y+����9�U>�D���Oe��O�_�/�;kP�2�f��Y1j�R�4��{��*A�"6���A��NST�U�_z��o�60�^��L[7c��ϲ}D���k��s#��R�$���Yg�ꋮL��\�?�xx��᫱�V�}��I鈈������F6�7y�^�J��kM�,�t���O�l�M��~v˒�Y���m�^�a2�砰Vݩ�����V�h�X���o�+�8��@�|c�Cc�O��ý�u
�ǗI�˟V�������XlPJU%6&�NC�SԜ#L`�CM'�䫫�e�^v�o�lE�K�U����7�����������'7���\o�L\��0�xT�X��	Emk=�>o��aF� K�Wf%��0?���@I�Q�Ԏ��ui��K�'[zRV�><Y$�Y-	��y��F�~�+#���C)���z.�UO��ۢG�u�D-��C��y�N9G����'������N�&��"Y˸�
��X3N��������TP�:�E�]�4fa��w.z�'�}7�;|���(���z0j�t�'�����Q�57ۿ�1Q�(��=��ף�Ұ_j��ʿ'#A�#�E�M��(�=�	��X-d[yB��u�̀�.c�Yn�����}����G�'��*�����C)�Ib�	�~�w��,�C'��;99W�%7����� 5� ���vO�o.%�!k�gT��m�iV����-U#�g���fԟ�ݟHZ����=2#[�l��Ì�k���d�����Rw]��R�"z�{�	�ǣ���h����b�kKζt��(����2���p�F^�H�v��=iA[5c�y1�Z\W���J}�ii4$(bSBGU��!MN�`�;�ݘ�(�8�ߤ��Y�G<��T�V��^�(��v��7k�\�s(m�H��횉���}.3�DV��M&'\G��DAA�J�a����#�ߝj��������(����6+�M���Dݧ9`6�Z�G��k'@!������]��Lѕ�������Sb[j��P1zJ��p�Ry�,>;�^����u* ���ҭșJ��Vv��(B�̚�J�����^����mHq�S���I�S�\1�.<������oW�D��T�/`bN^Y_�_�����AFB�뤐�:�N�Ý��l�X*�et�&s���_����NDPDtX�Ҫrze}���V%|d�F�����F�� ���]Ґ��lLvA1��]���h�F8@�
��%g��PX�,Rps���kw��\�M*�f�na|A�9�6Q1��`��������W��H<�/G�ႃvIb��;?�}�!e�vI�B��Hu��[��Y.���r�?L[�)K �W&H�J��5������h)c���n����>�����+���=V�UQ�7x&�n���P;p����ͩD9||��%YL�a�JS�@vLq�Z��<�5nj��EXZ�?3 #�L?̛W�~S�6�Z7y/.;��n9aqe���m�� ��|nF���;q�T@.o�("� Ըy8��R�a.󖯡͍ț+u?���xG�x=�A��f��͞i��ڋ����y`���1{%��&���@־��U�;Ly��z)q(����D��Ŏ=�_=�L�<w��J�ֿ�Y�`{c�=O�T���+�4���g�;u���Z����ʢ3��o%�z���\�ҿ�*5![�t�a�Gx'j��E��C>^E�M:S��/��5+�b�c��>�th.J�?Z8����tǺrUlK��}�U��/Ϧ�҈�\r���(�Y���m�罇_��*�Бsv^B%��~���E��J!p�D��y7H䓝����Rv�B=+!5e��E�~I���=�.w��Pw��RoV���w�XσxYPw0�n��Ҁ�\�=�ǐmێ�]ꐤX@P�͟��1dx�1�;�o���>(^��ޤZM���l��K�?H��L��Ծk�^x������	�����֟�^�	џR
���ҧ]XwO(L�oK=���f@2�|n��8Tx���h���@y*3Ko�����<|5*���qK���!��xpVH������M]3�sB͖:~��4C��.�M<�0�����m�J}-���� ϲ��Ƕ��]V�-&lΚ���J}��jr�6:�Pd#<[,��Nw�$,�ٮt4�������"�'o�?���5N7���_���F�V���ddf�$���#���"XWި��KQM����>ħ�X��<g���å�zo95��䎢�k�����
'L�J�6Տ4#
�ܷ%L�	���aU����}]��"Qe�\���x�$�>����,$A�?�0,B6g���+�v���q6�rVPCK��4OK5̺ە���o�FH�n'���
Ri�.f*��E2�i�߱t�p��}w̳�ޡ��Tǿ�d\��,�s0{��*���Av�w�Sx�=��ڻ�	S�����e}��U5Az��%Cg9�|T+��'�6�!�6�"��n���8�h��sR�G�ɫ=�αa)eԛ/�4�|��!?�m���S��~�J�Z_
���T;�
���Z\�Ѣ]�&ס3	�k�4KS:6��ZZ��n��� w���*�M��E��i�W�_�i��p�+f�eG�x�:�7~��Ս�L��F�_���;�`zE� v-�H�O����Z%6A
�e�N>��x�XPdU�D�W$۞�t$��ţ]B��ol�D��M�!}�R�WD����!�1�>�	@���W�����	��pY�u+�>!@��;�YH���d�s��"�C���c:�	 �Z(��I`~�o�L��p�Y�t���y���<auƚ�LkQ'�$���K�H���q�̝��NNEq��i�7�s�7�y�
罴/[�.<5�~����p{(�ْ3�AEQXm+��h�0t��p�%��&���g�Ɯ�n��z:����A�n��,���ND���s�U1��2%�ë�"��ʱ�縴��xw|���@�#e6�c��Ξ=ݻ�3�ځ�/\[?֧��|�kL�ZZ�t�8�>Z�
mu�?�ǌ����s
�1�ɰk�<$�$��L*o�@㻫J~B8�ε	?�/G��ȟ|`���3�7�9Y͹�{�{H~7�)S��E��H���4��HB�-����o�_4���U%*d��}B#´\��i�FQG�j;�뀹$�͛�f���ze���[���0o��Fw^�ٝ��M���)���ۉm&��2bee��%�Wu�}��O�B+1��>{�z�7#�XŻb�4���&w�B��Dy͜��(�6���ew�u^��<e)%�u"���iK�k嗩�[k�3�k�u��*�������"�W.�=��t�lL��Ƌ�(��%�BQ�'��1��l�2J���x����7�Γ�֝�fv��%��OGm�>��}��m��	OYk�}=��]	�gs�:B:���q^����x��T���:�M���Ç�[��&�����x1��y��7��K' 5�@�!�u'5��u� `S�����r�!Q4�ٮ�z���g��D�G޷],ѷ�����+�h�+W�:��ɩo������Ͻ%99XU�YҖ�x���5`�i���ϩ"���*b���Q�vǤs��t�L��@���'�w.l/�a��C�����MbX���x��g���� }kK�-H����0C��D{Վ9��������5�JtfCp~���vo��'j/K���t00�H�F�=DuR�U��\�*R��R���?��E��N��5o�[e���a�Q-�4�EW�(b�b�fՙF���8b��%��9�k8 �$�������N1���k(4bq#˪��=Z�W�m�1a�)������l�+��tUM�l.7���k/_�#⟽F���'�[�K�6�2"M��P�;۳n���8�~�bM �j�8���)���T�
��w���a��A.���b���������?�vw�{I��g�|��k%-8/#�ni���s�uH�ҁ��XX���Ե_���>2w�A��n2�>p�D��ǜy"A~�vX���w��Ч�d=���m{��w��C;A䵕�߂ǯ�����wx��GA�Q���g�u����s�@F�qy��!����.	���_+�|�	ը�������:
k!���
Lf�Ḝ�޷����`�ə*�ϡu!���@�`�P��ᆻ�p��B���u��"]��\A��0���盉��o���?�|Q{d45e�ǅ�_޿U�*^ӽ�р�W]kc@��pCg:f0W����#�NH��A�\�G����>�h��y��L�� ��<m̌���4�eM��sC�m�%���y,�M�OU	x�M���]��G�ez�`��8W��%��3�G��e�^�+sN&qR�7[�P0?,�.T|�����m��G�mr��v���q�m3�j�~�-��ѿ��P�y#�W�=*��[6�g�}��i`��L�E�kYV����X������<�[bd�.�-�ۼ3ѷӒ���8�������ԊlZp
�$1c�_���4!���Й�6�S߼�j�sR���A�BnA���l�W�dS����`Q$7�"���l�e�qy"�,��C�-���zs��x~���B}z�I��"j�'k[}�.Pp{Mx��I�s�ʫw�'߬v'�\����a"�2,�-:<���=-'��T@=h��%��8�s��l����ŋ�=A�Uv�}u����ەx��:���3����	/�D?[3��&1��Zt��Q�;4��F�i�E���.
v�' ��pR�k�9)/���5�c�,�t�i��∟E
�5�*xZ�f��Ԩ$��E=���$�Gع{ǿ�
�cB�U��u�� ���� ��B�ZC"��%����m���K���<�� ғ���ٝ
6f���W ���ܢ�W��^���>�َe�>�PK_Q��Z^
 4���ʭ7��p����'�j�m�CVb�N(ʼ�Թ��<�c���3,��g�Q{%�T�Ϫ�z٨���Q���h�{�=���[�И�b}�����U�#7^���ѐ��R�����ZCWsXA"ٓ���6������Q2�rO9v��e��l$����Ǚ�ɰYe���{luο��2WP�o]��F��<,�+�mĕ�s^_�Đ_b-(�m�a�����`9��z�-kM���Q��C;�{
{�	v+��VF��VS*'����(L)�60~���q�Ex�B���L+��OXΈ�y�?�+�F��_��
�������,`��y �a���(���Ulj�I��a*u4��eV���-�$t�y��ej|�f��L�n�2�eG?��K�pt+/�'�f&���/i�`
�Ȧ�V�0xr�휭��J��Ð���wFQ/�[��#ɣ�9߈���,�)(��yqE���I���t	���9�[�IVJ�Y[U������*�x���7�fϕ����描���_o��o{)5��h8wԓ�I���*��WF���)ߊ\��٪}�
6t���?�?�?��g�_V�lz��ݲ��--./:�ܯ�\����"�A�c��`-��ֻ��#��k��N�V=0>�6��2d�<w�CH-���b�"-EU�N�*�*n����U�67lSSV����/*~EKYL���e��u�͡�,�Q�|���~����/1�C};��,����M��v�����$���=�������aV����T��BV��S+G�HG�b�z��� TJ���?���[�X�3����76��l������~����o�]�'HC[�G�C���7l���^b�g\Ժ�c���k\7��� �&�á���01�~x��#uхȈ��H��!���t�q�h=����DJ�0����!�� t�p]�E lͿ���l����=�պ��"���@���i��/�H�[ޛ�xa�B�?�F�&U���s�9�a����ƲW9�`݇*9�*�IBʹ�W��O˙ͻ������ވ��t��5��Rq/m^";-]m�|���Xe1>Z}Tp2	�h�;�O+g9r̼1��Z���j�ZfK�� ��t�X��`&ܘ����a�d��?�)&L93)�h���̬�&�X5����#�Dq{'7�Wg��S��6H�ǰ*
;��/��!����[E'ܵ�*�|{0����p�ӥ��a�>�x�{��9�P�0��,L�uA"�|���T��t�=�V_5���� o�({!E9��~sj>jYԚ6�h�J�W�g���D9�"ߵ�������ڙ,�*ǶM��	�g8bܱujL�*9�P�� .�9�fs���R��.d���N�fi��`nl��)}ǟ!Ƕ������i���g�l�!V�,���:#�P����Ȯ�ڱ���Ɣ;!_�կ�p�ɶ��k�CONw���[�.:��œ�EV��]��ب���!����l�@, B������������	s5���"�L�w`,V�i�a�gg_ˣf�RzD���$�Qh.�]�����my��q�g؅����
��H��_Ɋ)��Zvg3��	N)��ο]�=�0a�[�~K��=&\�o{PWɺګ2�d�y��;&�������c����½}��VWxG��U$ެ�)\6'�>��j�6c.���i�n*˷�Yh��J/�٦B5��Ϟ(;|�mǁw�(Q^-t��6�]MdC8��Dx8I�w�[`���?�5G�*�k�'����iq��������$v�2u��I��[�n^��^��?Z\6��v3]:�#ފ���lU7�O��9�>�a\	��3�UK� �{RӔn���������l�N>6؎����.)�R�[��5�G��ni�`��rH��z�i�\`5��g8~�E�u����y�#2�R��5��9��6���8�z�u��u�>Rz7����.hV<����W�M�%�{���B4=Aۺ��ւm�Z(��=�^�>��"D奎׎���1Ҫ�@�P�X�y�g?F�ŨRh��k%����>Sv0#�I�37=�r�������݌��2��նȼ"�4\G]Ϲ���z:C|��W�Vc��U,O������%��N�j"�6�((���r�7X^|������
G��O,�_�<,q3�2iC�c��߀��<���ٲ��ƽ�-Y����mC���G"3r���a��2c��#Zus�h2����|�:��L(�j�'�M��)���Τ{���a�4'�� D��C��l��.Q���a i� 3Gr_�Q����Zd���^b������9�q%ah'��ʙ�B�^.���N��Hf*ԍť���:Cz���G���>ɯB�[cQ��Py���?���P)ѓ���'u��oK:���0~���)E��
�:'�=[��hd��@u4���}������5���g�}����^�a��TA-HX�%t�ƻh���56?�-2J�J����x4���T��_�F
��4��� c�q�_��.��*d�.��b�/L��2t��u˛̱h���D�p�qd�D&ϛ��f�&}b�o�Ą��| $����
�U�K�|��d�v��ٹd������;���׆�'o�:�Q�#��4Rc2H� ��z�%�Iŷ�YY�R����G��Ã�#x�Pk���C�����0{�/>���9�������5]�$�$_W��{;~�Ggqﾸ���hI�j�hD�̿�A���E�I����(�7�L�:}|�L�e�8Ѭ�3g�UY+������-����b�uz�_sb��;����γ� �X� ;Ҳ�/�M�W�_�*\2���ކ���~:n�����]Q�HY6?���O��>�����߉�v��-�7Q�x��¨�Z��Fՠ=�@=0�V
Z'Q%s7Օ��M��y�s�iI��x֭�Ev
+�3%8��ojKٹ6�xc,��K��cä����0����_rE_J처���h����L�Ir�i��z�V��j4k}�D��I��;��wbq��>�"�Ά��٨��4l�lb��M��9\Z�ɠ�l���Fh-�o��N6� �%��O�`Do���~�<�J-\?����(����ʉ��n��$��8�\��uK$�<��!c/�X<7)�/�<"^�y5k��g9�kgph�
����Gu*�8��j�ڶ�͹Y��T�H�5^j�K���*b�w�uf{o>�;��oN�jG�G��T�C\\f0�nxn�}�Ɏw)��o	Ox��M�I��u�r��>��k��6�N݊����&8?
�*8���<�C2J`�
{铰$,����]���H�ӡ�� �2-��o�!�?���H��;�I����ͨ�̴�'�;^��k���V��+��mZ�t3���/����t�� �E�R�K3f�j���_�I����c�7��եo"&�W���dx�A����۝��?���Qjrv�|��V[y�neW$6/�ˡ$5�?q٧rK?l$�����;��g�Vu�x����nd*�Mo��&��50�V`���l�jd�pHֱ��b�l�o��]&�����Lz��EEgPf�e�#/�t4DTAB��x
B��-�o@�7`ֳ'�B�Y!��7A��R��,9r�q�H��!���\�@�|D~���9v�Y]��t�]}.d�®z)/J�7��[�?%�>R�-�x�F87�}�X�k���~�0�����\���b���:A���|��2`X�hRh�N_q�BH"R�؇�0�,<r�wIr�kB���_��0��Z�]��d�6���=���	��|��2��p��rQ�-$��HS�	��� ��o��c�1`А9Q�4YH+�)Jr�ge$t�"��q���Z�y-�HUe�'�%��O�	�À6�1�tG���'u�V����>��\����ڰ���	�+���K��B��������EY����X����ZAQ����cТ%�Y���w֡ ���W�C��7�8%y��%�V�����MU�{��N�	��������$2�7����ޯ�,~�dC�歭��\�St(�Ҽ@umn��7�'t��_���|ˋ<B]���t������D�����&YF;��%����v��t����ш!I;��WNZ�������2E��9"mTkqf��R��2�'�'�����Z߹�����tp�\>��2�=��:��Z=�/��F���u��Q�k�GOQ��0�7�X֮)���F��܆�J��B��Ν-̎�sLY��Ug�W�$����X����c��Q���>�A��a6�����
�@m\�&�P/v*f`$y��"�
����5�_�lay=x�4�����1_o�����mư��9�1 �+m� ���[{Or��t����W2vX�g�jy��%�y�:�:���'-��p?14N[���*�F_�2����o���FZBJvӶ����<�	m����,��E�k=RBi��>Ү�6u�t���Y�1��a�ş~��M3��ID}�Ŝ���I>��U���%A��?�"���+5k�W81q[�����"_����nׁR{�H㻹`:	�@�Ѭ���o���W�j|�"eI>d'c��o}b���J��֨?���y�-���@g��t�3b�	z���ԡ-�/)I��QP������]�����`6�!9�����y�W7MG��r���"lZ��R�R��l�iVwbV�;炥���P�o��U;�&{>��cTtx�8JW��F�Cp_��& ���]����Ux�������Λ�	���b
қ��@����.>�m��y��8HJ_1%��/�k6l�2m�Ѧ�R︵��a�9�|�e�2f�G6�"b��������_�9�=��[�$K�zj��^9�M�T	l߿���K��9�b"��}[����|Y���#�pA"�A��9����|��@�T}�K��#"���Z);J�?JVT7�ػڢv��Ѐ��m��q��-Π'P��}�@K�Fŷ�rt�o�ļ�	��e{6�뷮�z�zշ[�ϳ�s�8��c�w6���q�Q���$��<�G�u��c�ѫ��!�>�.����O�|Ҙ��ә��{V���S,s��::˵�g7q�)`J_��Ħ�uO}�3��iyڜŇ)zde�%5�Y�A��u��M�j]$\ñ�4�����p}�Z/���7�w�x��)r�[����t>R������w2)_����W��� n:h4~��rV��=Aq����P�sz΁�~3����o�vCXu����v؄0�fjoKl׿w[�xm�"��EVJ�o�a`�	t!΅P��D�_Ώ{�*�B�=<s8�W�����7S���]�!S.�����S��f�BO�N���I�,Yaj��0wy���)g-@H���Wb��k��p�ˠ��#|*���ׯ-A�Tq�&�>�9����11C�i�ͨ�����Ϸ�)#Z��)D���v�y ���Z���~�J��K8��R�6��� ��f���s�FW@OB��9�T|P� P�1�Y��&]���e��̡�-?��5��Y�������E�}���<̍6$-��E��C�����<m���_@��t*���vB��qH�%:$���X���%���i�Ʈ��?!��c�~r��c�W!\H�2��#�mu4d^��L�=��wjXRùrJ�b��7I80�����"�]��S0�w��@����پ��>������3�Oг��8w�'b��;�j3�:��Z�9�A��4�Nх<zˈ�x<��)���Ue���p�!�����]I�� �p���x�(��Xo^����	ɴ�?T}w\�KЮ���#�DQDAAz�QzB�R�7�$�(�4B�&��^B	$�ޤ�J萄	I���w���ewg��y���}��䢛��[t�.N�I�Wx�gP�f��n@@�"�z�Ů.�wo�0����$�u+]��򛚣�Y��8Gbz������2������u�����kG��%}��m9w蚓��OЮ�E�w�������EG�-6�a�N�%�1�\)��q&˲ɕ�K��@�����Q�h����+���XǭL�H����`��뭔������cHO����e�%5�,��-}��1�i¢s�͉�;^o��L�Ӣ��׀e���\�#H�7'�z����ނ?�,����FMak�ҺD��~4iG9"M�A0aP�A�4{��]��i�X���Tg���.?����s���
*�X\��%ԎR�$s���U-��B���Ǳ���/���"7'�z�0��+��RL>�׹�s��.�)p��x��9-�h7FȑBZ��k�[�d5�MRG\������ˁ%. /m�0�Ï-�,ΠEN�wZ�oH5<����6͓T:?�:lé�Rc ��4�����7�}=�g��SV+��K^�L�n/��ϵ��{����=+G�������WR,ys��c�TuO�E,�r-e�����������q(";R��w{*�C��׽g���+	UQ&=�eĈ��fŦ��ύ�����_�������V�l���Q�-�p�̀d�pr�4�q͚�k<�N͗�2=h�t�g�~U����-eo���y_����fJ�q��	ǗU�������EM��ɼG5��I��dc����=�R3��Z�Jc��J�����u��%M@O�8��f�U@#γ�>�c6�ok��v�k�������x#�u�Aڨ�>�W\���FR\c:p��ä�W��"�s�ӝ�Q�Qd����HL f��@aw��"�1@��Ua���ʦ��&5�|�)~����"\�7�YC!�w}x������������w��9�v����I�[5C�җ8�|�T��K\tb ��}��cqhK��-\�dbF�Z�2$�&&}�u� 6Qw����'Ԅ�_h�
X#�>�٢��]�O�"ҸLM���O�����<���g��b����_�r��TI�.Ǡw��V�/U��<\�[#��T�Z��(��e����K�������ĵ8'©�g�ա�U*\�\m$�2%��`��0\��9�}��S�!���3F>�ss���sZ�@��Y�|�X@���A�����,@��e��g�������_mt��\5���2��'�ȏRof��fq4����4�������)֯�C������殹�{<�{�<6��N����y���ہML���>˷�cQ��0W���AY��|��O���m���>�!����d�#���x��E��d��|���ާ0e@�V[:�J�Y�P\��)�tg��?�՜�r�$��}p����.�)����L�J��K�!3e�lV�.�17D���:'�LJ������A[�t�r��s�b__��G$YǷ6�R�x�pݩ�<�7��V�Ռ�$%�R.q��*��X�_鴥m�;���#�ss�X�X�W���1u�o����A��r~{f!�Y�0]�����>7�,�#��c��(�o6�J�C�Zh�]��Ɍ~ڽ�~{ y�tR2{a�U��]{$�����[�I����Ľ�2.���:|���<�)7cb덀��ID��o���7߄W=*�B��6����6�jk����@�P�s?b��/��"�]e8���V�@��.�fb���W~%��3K�=��ɥ�I<���'w���l����O9īӆ�D�/��8�A+?��ҽ��h������3�'��-�|Q���q$��CEI�݅���l��&���f�@�O�9�}��_1�\c>_w=p��2�����4a����Uh���ެ�ƁNG Y�k]�^��rm��SA�_5�Q�actfdK53����A@t�6��</PC)�v4�,\`,=P�����hF�(R�3R���,�.|��X�<׽K:(4���)�K,H	��h�w�FB�V=����(��wVW�E��Ǣ ���U�X��L�����U5n�A�}D���俫h �����%���f��4�ݞ�o�M�l�*i�4c���5f ���aYK�iD���`���g�����*3y����KJ ���E�j��crײ��8��� tWA��*��;T�R9�yO�o��[�g��;�n������7T�b(o�{�p�,��n{׍����o	�R2���M�=���2���e M����2��y��Ƞ�7h7ˊMr�JҢwWO��j�vd���>� ]�L�i�N�|�]XYZ����8�J�)	7}�$a۞������\��p5����A��`��ӂ�\��^[ANv��	��0 � ��HM����?�`xz˞�_DB�H��u�
�{�'��+z+�c׵�H�O�4�2�;R{8.�5���~���}oy��kt}���$���uh�:i+��V�(�vxUQ��
���]Pbؿ
����H.M�5���D��4u���̴?u"-�M�C�1��7��OB�\B�a�21,�T��sb���U�y��d�7aҿB���ּ'.;�a����|��%&���\8YqD�/e���Kjl}�@~��^��>�h�p��D]n�;����#NdC�'9ޘ�l�w��J�.K/Z�1W����?����7�%R��Vۙ}]�����fs�sx�lLۣX�X�/-ߩ���֍J�-H��_��` <>D!2�3�v7�M����'�$v^Dn�g��iuA�h�e��8��Q��.8�u��`�~fo�ܿޅ�N�v��VN�;-�&�>pG��|�n�S�ʣ��8��#�遗��������f�֣s��яR��y�X�#-� �"a��@?��I>�?�_�XG��L�5��++/����y�n�����������ݷ��l��`�7����t?�l����J<���*���S:�.˫�=8���TԠ�}g�5��}�E���	^/BUT�N{�3rF�q�j��g����/��K]����Q]K��������歩Ƌ?y�b����ɥi��{VG�#�������P���;x�\��#`q���Ѻ�XLĹ����Ļ)�ӟ�;������}.�����~ ��G�-���$���芳�~�~�PD����2�ݩ/y	��9�Mh\_n���B:�T�f�8�P�]]�Ѭ��j����耕�i�.��7Ic��V����L�4�+}����Z����fR�L�z�Tۚ�q-�S��2w�"=j�`�y���zm`�aZ�ИF{(��`T��W�%�RK.I���9��]��Vóu{2��m>�n��\-ĥ13�R*ҿ�[�
��xY��O���ޭ�Em��If���	���*�i���y�� r��^�[`8�ʣf"�Z�~�}�[�"������w�����{��\x��ܖی����oFSK�����%q dQDAIH4����6�Ney��ӣnQ,"�l�罻z�Zfv�nMh1Y�Y�����E��/5p��>�+-<M BHk�_:�Qf�:��N����c�����7�7e�Fq���-Nƒ���w\��� �.�.�{D�, ���$�����˒�S=U~�#k�T\p+�M�["]��
�����+{��/��e)��R��\8]��J��C�QL�=l���U���#`x5�4�-���ҭ�fs~K�k��7h{�,f��bǡ��W�><ё���n��9,*W�)�7�`�W��X72�p��4�=�.-@`�I�&�J4�l��	9��k(\\5Il�^3�B�[)Z=襗.�����i	+��-�uJ����w%~(08�yq)���Ki����ѿ� �ɉ�����"g6�m,ID2>���7�|�6RYk"8%�Ĩ��X�y��n�oR��}�!����im����ǌ,��:�t��ٜ��3�W�ݒ;����S��s�4J�ٛ�L- ���]�v>��P��H��t*�.z+h�M�NG�Ub; �(Ƌ�xR��vl��rdZ�7RH��/ۏ%N~��($6wjT��@o���	��>�!�1���h!�Y��������A�:o��g���["�/�Kg�nM%v���fڵ�������׭	^�,+-:~�����{�ۃ�݌��	�i߇n0�7�8IN�G��OHG�z�4�aW�����1��i�;�y� �e�s��ۍ5��䠧z������`d���Ë`۵��_���s\얒J�V��2��U�J=0��OT;���ħa�~�Hx�_����7NA-������xN5zQ��+B�Y��OT��t�✵`̈���ߐuuVU��j�1�g�(>n�~�MP�n���]�K�L��aVz��]��%�/�q�޻'�G��5�� �e�6��rc�7��0X�Fmhl�%���I���������b���~������ɑ�9�U��^�v��q�N�O��*���(�]c�l����w��̬��6�,��T��lN��J�LM.���M3�ʕz��a\\]��Ъ?,#��[s<~D/����O��$�P`��6���I��`�?o�N�\��^���5�%m��[���bC�� 	��˫��w�:d�?��k�v�lv������@���J�R�lG_dQɑ����i�,F��%�2Bʏ�K���z������fd?@�'F�v��wB��-Y��q�SeK-E�r.KET��}H+3���'~_�X����!�~�i���yq��.�����I�F�G�V��狟{:ГU\��&�ν
#դ8�*�{��t���L&=�&	y��z<���e#�;���諾�o��8)���Xu�����$�m"t���A�Z�&�-/r5񥩽��S���"�5��tACG��Y������R�.��Bz��/�":μDPp�qH��c��1H��tؕ',��(M��l���}��rv������
�Ss�����^�O�u~�i��	u	���eD�i����r��wL䱰K��+^>s���������m����*�)�|��9��n&{zv���(���;���2���OF�@/��i|>��NP��-��4���C�ov�+&|
������u��ɲa��v���je0�F0������c6�{����5rr�Zv�z���[�.A+�ή��U�o�k������|�i$ {��!��Wջ"�	��b��M1��xl������떙!
�wõ�Kq(�؊>�S���e�A��K{sb]�d�����Wu�j�����B��#5 ���hr���9���v������x:%���{�>��i��Ƅ΄���h!�u��+�5�n�ć�b�;3"(�"z�k�[��6.l�Y�N�ąF67j���֤b�t:�6m;
qܦ����wY�v<.�#j*=�v>a*娣������+z����|��I�����uӏ�sEpћ�xl��وhȫ��CpP���K��fe�ɔ�k{�
�`b~��ܔ���V$��LfU.��*���bs���47�~cH�?�M�$(�-9��"t��W�Q!�ﴍ�-�����#�%,��\��������QTԴ0
	�f8Ua����8�:��R1[���o�&�gk� ��0bN��d�)�:�YvCsCJ�X�ٶ܆��	��.�����7t��A@,��k��d�.�I�&�t����e��/���$K�a0x���J�� �X8�Z�L�}��X�i$&MVb���Yg]�@��|V�TR^�k�[��j�Y��p��z�g�H�*	���_�h���RF�MvVm���%�~R0e7�0B�S�>^��3撧�Fx��i̛v���frw��Cl�&�y�{��N-�'��Ey<�X�G���%��㰺{R���f�`$�v���F�2#6e�|�6< C}�(ױDx����\�)�#�9Z*�E:d��>�o�:�B���P%2�3�%~�}u�o�K�N����3���iV`��U���	7�-��L�t5����04��w١pU����M8�-v�7���?��H��ڷ������D2�3�ҭ	��Z6>�ݼ�"\�N����=�/\�"���Y��@~��������lgsw��&h�7~�(�;���kp�{h�O��Ӎ�RDT����&�i���k1`ʷ����A��(�NNs��/�ٰ��N���e��#0ZS#[׀�6����Zh��my���7\�(��(�M�i�QP[Oq�2��GPs0�-rY(�C�o �5jd43Q��oǌ��";�%G��"��<�L���o��q�pŋ�w������̈'�����u#��iY��G�}�S��91㋱c)G�{qP~�%��T)E�e0�%���y�4pʢk�d��F�.��ڽ����&Y&%��B�2/,���N&çj��a2��h�c�P�ڙ\�a�E�}�X�<^��ۛ�L�a�b_ �8��b�;{�G/��/�i
��%���oE�.k�R�uiTNo9D�\�s2i|�B\kD��v�Df"K�~u��CĊ���Ы��*b=��v�iB�:���iv��kT�쬑��[�6"����Й����%�zٰřn�@��?M<�_��#9%~�*N��}���Bxzit�I��z+kM��h�7l��8���r�\�ȳo>$�J��L|�k9�(�A|[��>�f����VT�#�[��i#�/d�!F�2�b�|s:���מ�[5�Q���x���pt�1�ko�5�����K�O;睜8�5�
^�������U6>{����Q���0���,-��	R�5.�Kw���5��\�뫧'�u8��qq���vJ(_��xK��=�����G�q�t�����<6m"�%� ߟ��ǺT�2��9����w�;q�?�b�2`�!��{��8j���Gp��XsD�7�Guu�}�}7��A�y޲���ZA
2P�6p��1�X�)Z�-�~�޺���0�#H00���YI�V<�*�L75�\�����*W��"L��������v#��c�����@)x����䒟;(d�ڄ���K���S�[�mX7S�W�W��Z�s\Z}G�w������R�\ ԭ'>&ܘ�G�ď��'t䑳+7�Ւ��I�A�2 =g�z�꩚D���{۾~M�h�G�{���+�����Z\61��V�}?!G#��b��oh�gx�����a����UL�yE�R�{��9�\L���%`XW'����lR׎@��E���EQ����sPǌ�MQ�XGb��������L������'��+�4�6��r����uV:V�{;�s�6�в�	���fJe��1�޾�9?l�o�w�\d����e� �ʌI��u5io��8~���~^o���m�� �80�[�S�66�d�{�Q�bV�ublO�z��S`3�6�2gxS�6��0xP�u��V~����(/8'M	2�N2���?��^��g��]t�
� -��9�L�N�6�9��Pw�Y�+�!��~*�3Z�p:���Y��^��Y:��;:�ƴZo^�[)�`0�.�Y�����:(�>���I�������<g����]r�7ݴfF �FZlb
�μm�J��h�5�wt{�V�BQ��ݍ4�v����e����h��>{�q��>���DTPC^��U����n-�ɻ����4\�<gN��u�	ܩ�f�:q� ��c)��7��1/�r�����e�v�h�"W�+}�~�fh��1�Q��b�gt�r�m40'���9���Pw���O"�O��Z���"$���o�$tq掆�j<a���6����ۖ��_�eX�U�J�����p�����3泇Wl�����eڦ1����Y٨����x�M��\�a:��ƨ�:ܐ��;Ca:'�.���l)J�j?rI1.q�F��6�"=z��@�ٯ��	�hٖ16EZ�St��M�_ e�6�'b�4p�-%�,aR/�{�J>R�߲�5"�7\���I��̬w'>��nEJ�c#��8x�(S֊8�c�0B5=\NLl'9N�ת���
	� �\��z��g�ʚ6��.�I�����E �ӟ}����f�w����93������i�W)Z�m���x/�~����Kfʡ�kH�e�|�sjhh������;���h���լŮ	٣�.除�Ĳ����Jg�SRgz+SsR"����\�D��KK���|̄�C��2�ɚ6��3~�տ�t�L7M��_hh�4��֮�Ha&��x]�CQ�#�ޏ,k6S@�����Q�0�S8#�c�*��������vz�g�Gu�D���A�l�|}D���%'ˣ�#6U�����R�	���Q�.��&wܰ��2q|��kb��k�I#��-�;%�](~B.�c���.�����*�<e�����@��d�lxS8R�<9s7�nvp��]�H|B�r�vz�j�� ߟ�����kc_8*�s�$��3�1�E�.�=�ߖ&̵;#���p���0C��gD�����~��dޮH%�#V��)���y+4q�&�r��B�N�y��j���v�*�>�{�s�l��uԮ1���ߟu���I�
�� 9�ۋߚ4�ۣ�:�7�o�?���� ��� ���*�.�%Zɛ����2��V~7]3����>5����a�^�Y_��j���������������{�QOm���3Q���̫���''`^--�1C����C��|;�1A5mgO�(M�7�E-��JF|Я�̳Z���l6�d�	&m�[��we잓A�*�뫋�~'cI���f��Q�p�CɄ+ �Y�S��~��>��ׅ5ؽ��K�X�u��ΧR���"���#C���]�m�����)�%$����
�P)�?YY��	����b�"�m�_�G�GǏ{�s_g��j�{�G����s�2Y��78A0L�Q�5���� ���K-0�M�~*(���&��m)>��߲ �" ��R�%���-�k�`�p{�?/X��)$������T���5�c~�@�8��#R������V���Z���*n�����kÞ��������o+ܞ��	�?���f��hO ���������J��[��ϑ���R��M^
��
�Cu�Cd^���/&Īf1�K�[�y�� 6L_�Q�����R��
��1����VwS+��<1LFV�{8�}<F�����+���j����k�ܪ��M_D3�a���r���
NL-��U�,�؟ܗMa{���fS�5W�uƝ�U���(�<�h�LCd��xˎ�_5��`���D����̍��>p�h�� ��RI@�I�InD|�,?M���)F�wz��GT5�>�{��{��6�[pd�G_�R�G��̊��֟��/2)��6���D���K�M��w�����O�C��T�j��yc��s�diX� ����SYT_�&���X8v#>�6r�*�#oee���q%��f|i:j��$�⭪K_F�$� ���h��n��S����҅�^��ݍ=ٱ́E�A��q����z��Fy��d�UE!n0)*�L�I��D�*	��ŮaU�z�*#��}�zu	5��NG�yJ�(J�D4��S��E�?|��f[�{r�E6�����y�?<�!#P׼�
��=��>��`d/�	~w����VZy� $�2���c �Kӿ\���HH��ϨT���\���B�ڲ��<SƷ�%Ζ
	&/�_م�����KΈ�=���D�ǖ�xo;{ڈ����M��T	�"�7'�?�wz<��"Ɍ��X'6����G�|d��;}�q-Ɯ�a�w��k5y�6ܲ��A���Ûi�	1�)��5��)�IÔ�J��I�N�s=#x*�،���ɝ>�׌}j։��һ듦U�{[#Ԯ�D�)�I;O��R0�o��P(�8��+QH�ڦ*+1���a�޲���6WD�nWO���C�>Qf
�ߓ�3��������/
4'򹀌�Ҫ�h��?$�!�N�꺏.��KxC�n��W�M�R6��D�y>�|��Fj�R+��Sz�4��AH~���B����-t�<�=ۑ�1{��/�C̔t�(�F�ɿ��|{9Nz$����1OtoG�2n8�/���ڞ_�r �y1�|�:�UK�ZXW���Zo�N0c��l�əVg����|�����L8����L�#�k����S����W�G=��r�eJK_&�H�W��B3�F�;1>��o6��śڤ����Ό����'�����������7]�9.=&�r�K0���Q�B'��k��f/��Ӟ�)[*��p�8;S�Գ#�o�p/�x)����C�# :��5��}��|g���)�3m�A��5akp`"`*���i�T���a� �Oh�����n�$�+Ԅ�B�ix;��8���O����'��{،X��D�o���s�n'F�B���Kv�k뢟/��V�E78}�&s􋋓ʓ>H-*P�p�.�锄H��6���E�&�ۦ���AN1���>���Sc���dK�e���x������]�NG� ��^{l�N�!�v5%>�#�>ɍ���S"G0ۈ�^.υ�U�,ߐ��Ti��30Q�E� ��ef.&R�, ��u�ug@]gFN����5������*"�:�^z|5�D�DԿ��S
��|�R�F��{�dV��d����S�ƪ���5a.S�R��=�����d.�5|x�jݳ�=.qݗT����H���a��\#B�E��Z'��q�nM�
�2{�����ƪH������0�=�F���d� ��DD��؝>!;0�1eդ�+b������E^���ˠ���q篴vڤ�$�>������ǟ*ī����`aM�����c7�2������E̒�����x��햰E�X��z7������0;CY�_���rر}~�"]�-3�_����\�,\��~~���גv���Ǒa-#��H��B�a�~����h�m$��3�å��&̷VvhݶZ�,�FnO5�=݁�W���6фP;	�u�O�S!�#��ƎӼ�~��hHٽ8���F��I�����~d���'j�0�$�13�V0Գh�ա�@\ATDMT��ad��uflgn�#��l
ﰹ�,��w�C|��<��N�_����s�0����k.�;F��EOo�$T0��*�=K�����Rm�-�;a���x�F�9��3MΣi#8���\3I&��-�J� �դ��)\'���!7�"��j�k�����yR]d�JI���tf^p1
xw���\�LzhK�צ�=�w��éտ�٬X��	���,���c�J��*��jr����������#�^l�M����ɋ�%b8�-����Y���U�xVo�ho1�����*��HZ�s�F悼��$k�O~���|hg:
�y3�^��:���ώ���K\���g찡f����W��-VT6�\pޝ��gl���{�:F� >^K��o����wV=����E<jy+{2��EMK�ˬ��	�o$9�bF�,�F�>I�oe�,k�Jo���]-����&��+vu9�����6DP7�n]4u����&��*�o���:�5���_�LRpNY7~�ua�W�I��3�O�r���H�ٌ���Lp���?�ƺ�_�����
աBT��\��*dE�"��7@@B�ű�C���Z����7�L����P�,��L��G���M2 ���������[� �n��0����V7a�)$��Z:Uy�>���)��`L�� ����~_wx��R���D M���v�
���s��3O�ht�l�����v���g�3�g�9��e!��g�{y��t�n���Y[�9ҹ���Ժ�% ��>��ybް�w^�9s�X=?����@�~Y�ߟƾh�='D���H��EK\Ƽ��|51ܾ]�L`J���c�S�`�ֈ8�m�(�ac)*V`]^����+��౽.;nV�OcX����Iqx��N	��'��v����A���Ԡ?�~��دsK�u��-hK�k��iR^��5�(k}T4C1,��>0YuV�]����v#E���{��DV�ؿ�IwVf߽�ͅ/R\���ʲ���7�p�d�K1�Y�����#"��%�L���J�柣�#.�~��2�dCl��Q��KD�/�!\�ê;>��f�H��h��P�g�!y�a���]�W�|�!m�](M	����Ϣ�g��1׉�K�&��!��<#��.��&q��݈oB��5o!�x@���v�EU+�;�<X�c�����N��{cj����A�� ��nD`��C������X����<��n鋷�56��4@�ƨR0���;k3?��B1W��M���x�;�q�ݒ�X�A����\��'�R:օ��䆽
��̏�|?��WUK2��]Hl��wN<���<"���eK��K=˝��5mf_"�\����k9�9��}Gq�>�~�:�5�%0��iBjvt�����R�eդ�9�����f|{������lt^�~�_�q��T%��۷/ˎ��۬��{虰���:�B{c��m�SI��
��t�3oA6������-�ϸ��ֻ�=E��G�W�c�︹=W=��Q�>�<��T�����}�-���,���>a���W�����B�*�!I?�s�hU���a^�����+�VyM9��yof��d���^�� �+�����:�]�͏�eGs&����E���np/���.�����:��q�Oc;->5H2e)��N�5�*¸���/S��c#� 4 c�J#lo���A��A�_������������B�ʱ4C����L۝p���:�Ru�&��P����&�@�����Mo��^o�}&�ZhE��^O�R��K�$>�zeHi��ack�07$�̐F�ᕜ**kx�.�/ 1�?� ��=����^��ɡ?�7)���mݵ�C�kџ%|㒯��}���^�`(�z���aU0�̆��:�{���<�c�`��h̡KoOF*ݒ�1�6ڲsh����GM����]UQ����M���j��C?��'A��L�.�m_�$��:��o�$�Mb����ϵ,9���c�]wYX���x���[sU�up]�5J�.��ڲ�G�ᅾ�BGׅ�:N�\��5�������$���'��//d3�td��r����"�Z��Z���[���m3�r���,Qh0��y�ЅӼ:�(ٰwwD���R(���+�_h�C�.��?t��������������-˵��X51�ޤXu{f�>w�q�iC���w��5��U#!w�QW�0M	F�!p��>z�'ة��XmdJnfV�lnB7'���,��Ϗ�f1��hT)`� }-��Y�ٝ�S�jOz�BH܆����m���o��Z?,K�[K��\�Xl��D�S^��6q�U�r�=��7�-����nR��ZS�Ꝋ��1�R����,j�i�x�S:
��%��d��.�zr�S��B��F�1�7���[Gl��8GXk�L��;���/g\y��^%�"+=��A�NF!R9:���|��=���k�X���#�gϑ��=^�	;(P��!zs�8�ߕ���NY�mY��L����z%��d?4�ƻ9���a%N	�/�`(�[����&��V�)άɩ������ŝA��`2Hi�Z�����Q��:ѩ�v�?�x���H�ϡϽ6���*���D'I����v�$]Q�����s��	�]�~mH�D;�78P�F���|�w�6+^Xo�	��5�*^T4�wz�\�p���/��",�@��c��b9,#Ez�lj{N��3�_�!��y���Z��^T魌�0� ��I�U~�ʱT�qcVk���͞� ��z���H8����_g�{#��ٴ^�oQ3e�*�maI�%0J������9�v�����)��ו���̎�Bp����c��; �`��'��M}�y����O���{�
Ń�'�����Gv<W�d��S=7��	6�H��K�/��@w_��L��c��u������[O�X�c�~aC7VC��
'��̥�^������[7�Q�(5ƻ�s��/廱R�����N�{��3���׎��$��B�N�]���F�z����KuI�Vtt)�\I&���6�0x���i,=���GV	�y��ߎFho�Y��(6�N6^�/�{��d�چ1�0����&:�߶XWc��7�{G���%��ko��p9T��O���X{���~�M<e��(u�ȕ\����%:{K��:$� Z���}��/s�{?�ɗ���(�y���� ��wk�gg��ox����N�g�Wӿh���rWjc�k)�<�id>ѩg���^����)W��m���/�B�i^Dۢ�Q�n;g�?�?v�gK�jBwj�3j9w@14p��:�pf5�Xx�]��S ���N�h�9���4\��V���@n0|4�n��up	Xi�Y�o�(Q�Kؐ�5��y�5�*S��)��	��=b�)q��B��� �����F)����M�1��-$��z5vd�\���d,�Wl~�'�7��� �:s�%B����?U�YǸ*#�I�f^�{)�/B0��K}�v9_V���sn<'8�l��%����|{3Pkސp�N������������r��::6L�O
_��?�C5<Rح�X�Ȝi�0 j�G����Ĭ���l�9�VL	�t�Ww��n�����	��5����'�F- �!u�;
��?ah͔��P����CQ,�ؙ׳�;�ѻ*�S��0>��]��ՠ{�T�+�;�}�Un,�LM��2'�K�����
(��L����]B%���Q��E��ٟ/��e+�\� �k=�iE�^��R)�qT�v�1X����8�����.����q�厯�ܝ��1���`�t���h�Adxs��rl�'���׬�Oo�#���]�fQO�u	�]�b,��꒶b�Me�~*��?O�ܜ�s �T�>��]���
��_U��3�Y���|�k���#�/z7�9� E�����R �Q_���@/�fE�"~n��0sR��^zQ��z������4�YR��Hиj����Z�W�����4��V��{)%ѝ�O0/�3y�A9�Jxy�n�״%����J���AS^v�P���w��j6�U�N6����*��/շ��c��_��'dK���퐫2�&�8�y��I�����?���-���mg�U������ң��p�ȝ�)�1N�Gּ�+�j�;��&^�wW/�G�e���o�|��4@�F��[,.��𗸤Oz�/�Os�C�Y����Z��r9j,dY�p8�'�k��;���H��H����$��^�ţ�S��l�:� {'v��<���jK�[1���2/h�}uͷ-��'�/G�oK�Ĥ�-���͒����U#�'�yyG�'�Z����^�q����M�N;G_����\��jCl�K�|�Ri�
�����y|.c�'��8�M{h _^�TZ�݆F���N��<�l��	W��r��	���vk[�u�O��&x��I&���uZ������<�r�H�D�e��qGq��c��J����w��{�b��i�&᫪�E6�Z�����u�K�fa���m��bæ�ł�1���u������Og�2"�~Sa�n�>�#�K�d�QL�@�;j`��[���T�x���<�nӯ���«��}��5�h����+�����l�Vn�0�5m�G�jw+�D��E7�/h�/Q�ʹ������#&g�(����釒�5��H��`2�C�z�_�;�AC�\��9ѬY���Ѡ�y%ɥu�3�7l��냯�������e1�X���`"D����4���1!���S�'/�'z��7Mj��5s�+�z> �y�{��ݹ�;�BB��*�Ȁ�vXΪX�#?3�A���Q�݊w�:~j:Z��;IW��ƫ��{��/�7n���ּMr�#ĂezK�bٱ��\�x��L�A�=�/��©-�H��y�_V�/��kyb�F��2��rj8�5�ve{l8���PK�)�cެ����r��(~�r����b?w+p�S�~�)����Z��O���y���v��7��Iҿu�O��aH��G-�t�#��U�鱈+{���rO�/��;6���5b]Yw����M��<�Q5����p�~��J�$wa��ãD�{��SPg��F�|k�;)����w�V���o�5���8���*ì������ve��3#xw�~I��1U������~��\���dG�}d���?*�<Y���P�W\@,�a�?_J�B*1�lem�%jt��.�3��%��G_�j�����lD��>N8���t�2�W>�_~��w����g9+jtT����{s���;,�u�&�|YJ�����C�k����F>�Tj��|��̍�s(�t����L��i��V�z��=�l��a�=�N���]�Z�"���R�I��k@�=!@�
�H  ��I��^��=�&��������*�f�3s��sϜ�$���ʑ�&N��,��|w.�Z�j����7�w�Y��l�-S��"K<�z�k��ȀPu�*�^?T��h�C�..�&�,�\��sFi�;d���k����a���N�K��"���R	�b������Dު�x]���Մ�_df��s�c�E��cI�{P��i�ּ�~�b�a��^W9X��=L���:d��0�}1�G��+��ۏ��`^�p)����0��9�G�%�'�y�V߅�\U�Ff-��(��/�h���f�5��F/k{k�%w���#�օmV����.��L� �{"|6Ϩ�s��އ�c�ˑu�p�vи�Zxrw�����sj?�6�ƴXy�(j�[�=
-P��z��"�����{N�����߮(��糇�MZR�%k���j�*|^��^�C?Owa�͂���ä����.\2�+[��+(���)V�֨a��HK�5�,��_���զ�h�����jpHl�+U�A"�=7�ۻl��y�_�N�gb?W���&BCW�^�[�0��.������`�K����n�B�q�Q���2��ޫ�_�䥱��
}���>=a�sk(���͂�Y-�i��Q���cSJ�M�Z��DXg�o0�TmN.�:��;qq�3�yi�r�>`W��|s��H���:@�����9�b�]�r��V�ua�E]�'�`��V��t51e+D�{���8�
����I��Ӳk�I��Q�A�zt�s��(愺Ԭ	�@.�nC���p����i���$K�l/��h7Ot���^`�@�^�|/�m+�٥�U�I���C�p��a"j�Յ��ϲ�H����������Qv����u�-�eC?�Rd��tl�ĥ8o7�@Mqeg (ҍ��%��4�������*3��ʮ].?�0��K+'��E�L��?�/�F
w&�Ot�]MX�(}ӻJ$��\��P�:��]d��ڊ�4��p�9T�>�@#�ܸa���!��}h=�Oջ.t)[��9���ձD������[)�P�P4���2B�g�Pg i��v�Ԯ����c���rʶ͓uֆ8q`��Q��uѥ֥^O��iٮ���;�'f�fuU##��s�.���4�S jS��Ō�3x�D��X���4D�.�W����x ��V�{C��*��m`����ԅ8�c, ��y3�u3�LS���&�*��I8V�%6cS%p������ч�BaNl"\��)p��4.L�٬��@��ʗ��O�zor҂��C�~��f#��_��p�j��^�jGQ�-Rh���C�R������U�댑/�J�mC���K�iI�Y���֥`�|���s��V�6C]@\=��T��F�$a�5�A�=FU�-I^����n�υ/'����Jq�9k�4B�^KƵ�a_��Ԉ����dI.�؅ �)���>m�����o_�7\y��F�� �i�_���^��e/V=����a�Ƽ��Гp!�WL
|��l�����p;�0�UՏ/m���bR:͟�ؠ����!ySהnǝ�������o�՝���Y6����7� AR��ʞ)ss���O��d#�˥N\����n�)����|K��
\cW(6�3tx��׈���͹��l|��;�Y����!:$�7#u��gM҇��;��*�ps�D���D:Z~T{���C��$��CW�羪����|H���3������Y��<�X����Ԕ��Uj:��G��{�х�����ø�
��K
���V[hE�b��
�!pE� �}(x��黜��e�D�����Я�&�\��W��)��"J^������d���}��dEY�v��rR�i�4xˏ#ib�<Q�F��0���0!��l	ռ�:�n�C����d�s�&��)R�K�1CE�=�[D�280i�kŦJiv-#����o��i���C���?�w$,{j'�e�M��>���[��������,�W��3X���ğ�e.H�޽��F�ɹn�*��Ș4/1)���8���ܤ�׿hFG�:Gu�W�b�n�ý��[5���
	�F5:S-��-�Mή5s�D�x��8�"�Szkm��..�R�O�P�Ip`����wkƭ�0��y��y�C�Fэ�#��3�MkҿЈ1�X����W6T}R��#5����t17x�@���L�+%x+V�vp��d]~��u�M�U%�]�T�y4ݏ
�a����.� Di?(�g1����z�ق
C���Z!˯(�WK�ϊ6�J:N��'�<�:_O�5�R��^A��3���W��0��-�WIT�s}��_2(�gR�3���
��$ۚ6��K�G�&q����WG����c�=/"Jjj��$]Q<A�L!���҈�������F��?_Dq0Q��C�>���?n7�e�Iȫu�~����2����_�1M����u�
%0��@��o�f�eJgB@�IuY�"�q�����O�]�װ��ݯ1H4i��u��ZKX>EX�˦���.?֥%�%~�h������]���8ȰJ�����:�(Dp߹kE��-���>;X��?G�W���ޱ�41���M�s.��j�zz���ŨM\�� t�F��z�u"�Fyr	��$���oA�9=��b�ԓ`W��2!�eD|T��"�n� 5H�9�,Qͽ�}���>سr�1�#�R�����I�<5cE�4.���"B���.ўL�s��@X��	���̠ζ�J=�k�������axű���Ǒ�R.߰F������4!�B����|�a�N�^�M���#e�Y�	�p���^?La��������h���l�A�Hb�1<��������j0<C�ꠓ8����ˋ�߇�3w��F��~J���<\���ǁ�{�����k���M�����~;nF_{��~Xb��jV)0:���$t�h,�K�"mӱ�����J{��� �z�)	!�͏M���]�y!w#mX@CF�_�A�}���Ϸ`�����+��l��ZJ���C�z���94�~��!�W0r����#�=z��2za
�
�3��?�5$B��t��Y %!^�%o� @�E7"V��r2���r:���;�_0Л.�1���*w'=���l�� ޼�қG5/U��g�/Sjt�s��`Y���E^��/�r>;�pwmC�UH	�z�<;�� }�Z��7�p�|ol�۳W����g�:%�����'}X@�m�o���E�9kE���R����9�/�
�AOE�W��g 1�R<��#v�p��9��1-�9�͖���"�>�r��Y��=�覂i��(�Y��a���L���wFz�r�E ��Ԛ��Hw,G�^j]1̵N��� ������G6Y��.8Q����@�� ��G������5|�1>�kIl*�#Ql�hG�D����qc������}��x�9�K,4�Wp���rG�����F)y��]1���Y�T�Jw�oa��p���̉:�1��S&��R��q{��ļ�����{,�*X�Q�?�������y����@7����$�?C&��Ǌ��(O$~~��� ���[m�)<ˣ���#נ��8��3���
�L��"H��$�P���_�u��������h��IT"M�g��n�y�
���!�Wx�����nu�WMƵ���g-���p����#qi��ǫmK�.XQ�Z�?聜<�`��t���D�и��s��e�<���O𫬈opӑ�:)_�Y�%ʢ�K�h\�d�*� ���z1#��Rqհ��p�ɠ�]@J3�$)�Z���x���=�m+�7����0Xx�t��@k�i��c*!�I}&%���
#Ճ�ˑ/��ת{��k��=�UT~3�}>Y�b��pA�� ��GX/BF䑊;��W(��V�����g��"��vy����/����1�����G�RSa�.�<�Y��z��\S����NA{�+� ������<^���P��JA�Q��)]���D=Fb�)4uy��zx��i�������[���h���M��\��0���I��I^#n2��'�Y�g�=x�_��e�yyG����XJv|���4��Ev�맟y��Kuab|�=�ZP�Vs{�V����lm�����(:���'u�4�/?F���W�r���� �X�C�-+� ɘ>�3ô��U�s�W���az��nܸa>�!�{U,ϩ�9O�
����@Z���J���Sk�z��XdB�lf�4e�+ۃ���Q����Xy\�TP^�V�%:����C��)���0n!k�S$����×�"3�O;����v3�7�Z�0ZۼvG�2�"�(��Z���;�a5�SxВ�s�~��Sr`���-?D�b�u��܉�wdU�/�8,C^�rN�r��G9;g͟Sk���&:\�v�>;˵���]�z�~�CGm�B��j
ԭ�W��ʧ�Y�=��y����k������f}ѪH���Fraي�"N�=HΤ��&��3s ��yW����˕����ot�:�9�-)۴G���b�/<�y��Y�]v�h�<-t�'�:�>���+𩁢:��#W�
x6�i~t�|w�\���Kk��pgke}�Ɨ�=�pZ��q�As#)�d,�d���C
w9_��AQg����ƫ��������O<g�Ѥ�N�]�+�nM�Q\�����r%E��|����Ǩ ��e����U��R����v��zZ*����>m>�G�j��a�(O6���Q�s�}7�0I��'�ݶې�°`�@ųXf�{������Ub!�kS�\Vu�G�8K$�OY
'9���s\�"=���o[�j��S�J��[)�������"��龒`l������K��C�����ڈ���BP���!��8�؋�nuy�Y;�(��2d|�n���$C,#�l	�M�┳i�zI��s�>R�V��֜_3^.=�of�8�P/��)�k� �R��̷��X(*�7�z�E�;i�7c��d���M
�2𜆈k,˫'Z�U& j��Nˋ�U�OPft���R{翑��%R4�*=XӮͷ��@��Dv�􁔢�z1�F�Yjg���&�ݓ���tr²�JG���=��l7�z^��z��y߇�)2�1��;zso���唛Lz���J׮|��9�V~�r�t+v3�1fm>p�$�\���u�qκQA�D�~�MN�qH�k�_g4!��������w������g�ciS�X?���_�fwQ��a���T���Zr��l��-J��7�Bu����|����S�)J����E��9����R�CÒJ�Ep�����T�'!Z>E���6�@[���q������O5E�op��ݪ�Y� ��
�Sy����3�w��d5%��/�5���o�(D��C�W�"�hFèc�f��&RH-60傑mh���)$���Yۗ
��cu5cEk_���
�8�p×^u�.uS�(�qF���nL�����"�wȋ%�Qr1������=��J�)�Ù����h�&��g�]�����{#�(�ې��	�<GM�[�E����z�/��}eb�G �_�h�2<���`؂C�2���$)��!L��lf5�U�]�Pi��	��ޜ^���P��f�r�&VFG�$����kc�T2 n���-�'[�$�F<EhoE3k#�.}�-1?W�({a+��a���\�c��W�!}#n���-_/$f�f��?�G�J$�K�G-ި�Y��6!��Tr�huR�no���kjJN������(���$ �����_e��$��뙱��D/Q��@4��L9��:�sP*zW$�"N`�Ԧ���x�L��u!��)�����#N�STn��aMb_*p$� ���;4�&6��g�V"i��j�bkVD���K��YE������%,߆�a�#�ѱ	#�p_M��t �w3��i��޿�9 }�
��i^�c�&��-l��VJ��I��t����P\���]r"������xe��o�4�P������?㩎:��y���͜mr3�s�̨�U�k%�y2h��i��w�"�����<�6�~Itw� ���GN]K��;^ ��Rm�>�dF���K|�����%����m�F��G*��/8���85xg�It��v�J��)85�{F�"�VR�%p1'OԸ��g����&���`��nO�A�D�
(���Z9�l�1w�{ �H��0�� �ݠ������½��F���}��J����k[��x�j� .)�*!qf����*�x	<W[广G���&�[��'%��+���q��qI�-w��iG�!�dv�o51�/M���h_���3v+՗�D'&�J*�&w��ms[�ǡA��"��]-��P
kz��mj���d���[��z�;i{ݝ⽇(�#ha�CX.1�s�; ��3���/O�V�����E�UNt��k�WR���U*i���b%n{$m�g��K0$�fm���My��,AcJ��IF<�;��0�IvVh�TBuV�4��v/Q��}�[��v���=��E�f@�n{�7�m V��-���0��@�i�C��H]p�у����W�/��.�����D3%�1~)�� �<ڦ�%���@���x��t��T*1�y}����Ow�)��k;7�Y�O�^��za�v���犆���7��??���d �9]E*@E����=b�	��A(Qh��JpJr}m�̞���^$�~��)��^c��<�!���F~5���p���1�$�Te��``e[C`h��ъ=>;�(§�E43�9��^�B'�xq+�x��6%'�����er�y�����[LxߙM7Fם�(�C*,�G����|�j�9|-mϑ¢��HZq3�Y���\@�|�&+
fu�D��>����.���e� �ѧ?����y�� ~�Og�ժV���;b��3�f;G��v9`��)�@�đX�J�DJ/�����(���$,�t����=��31o:�w��yWaQ��l������؜��5V���G������B�m�;��Al��ڋ���P�qP�m�Y�������r��F����^m�n����.v�U��n���g�Tt����K{��qr`��t���AL����2�؅�Z;��d�+6n5��u ��_j��6���h�/�v+e��5��2��7���ǷD���[�a�|�7�G�F�%��[v�'멲�nuo0¡�][��d����^*$xp
m��1*3�
�H9����rOgGl��Q�5���X�_֤v-to�3mJҥ<���<Y�����2�O�a=���Om�a���u�.7��y!C�*v5���v�d��[􈘰/Û>&x$r�D��U��-#���H�*�6`Rq��烈X1��^�\�b6&jBob��F�Ġ�Lg͌��S�j?��_��<	���ZI�!��#Թ/�\�N�4=���.�����!�ة��V�o�:��k5�l2��[{m��&��d
�W�h�=�&طtx�
_���#&??�$���!��P1��^��91?c(?a�{�ymO�b�E%���Q�y�I�N9Q�mf�$�`y�i|-Hc%ϑ���T�S'�G��NU�ZA��f��a]�1z��(�Ԁ�M��=*�l�R4��5ܺEO��_�Q�OK~\�V��5�N���桳����g��O~6X�W����B���	0�f�Eabm��'�� ��w�$�B�Ψޔg��|)��)�~l�@��ų�ݞͦ4��6&}�ͫzDf#A��t��^�A'�iMMaK��B>���lG�;�����v��7���ۗ^�~�-�딦��<=�ᾚ���U�`A�=�@�R�(������IЂ�Q��4t#ì���m��*%߾�����{����m�}�����Q�^��kI�֝���{��d�k�w�܍�)�p���bAF�I�� ����kT�F���΍��QSz�#C��u)��x�}[&���,ҿ_n�c�
�Y���PǤ��nK.���t���j�i�(���YYE$H�ﯮ5��H9�e���ǩ3��X-e�F!{T���Rt0��f��]��e2M����K�g��4��<�d]˽~�O�����7K�C��PDk�"q36������@�_�{7��W`PȟFg@�olM�>_��/�H���f��!�������ޛ��S�aHK���.�ܖ�Q���T��y��?�]�����7��[PN�ò�B����� �"c�;&��B8��bO��k���|�`l����/U��^Eu��}ʄ�8m�	��>"��sR1�_�	óEwf��W��!����5����B{Σ�/^�M�;Jc/���Ҧ݋�CT��$T�8��لZ�[B�ʺ���rt���(���y�!�y��f��z>G��̖E9�;��sX�$�a�;�]0��K0�ޤ��$��p}����]�=����&��9\\�1j�]�����4V�~����l��4C�y-+'��n����]�?�i��jh��Fk^��	��P��B�\��*�<�Lo�������b�{T�.I�%Ϝ�����S:�K}�L9�N�/~�d��	�'xT���[��zj4DD�X�	���ey���u
��(#ۅ�y���S��^�ч���x���z�WM���vh՟��~lt^*3�,�eo�2!~���'��GhZ��_�����6�R�ʉ��i��OZ�%���*��W�a*�c#�@.��_�<�<�כ���nAvL������]���l�d2��h��U��R�������]�g�8�Y�UP�V�����X���%I�����E��S?N%aK�ҠӀ����m/Y�u�<Q4e����tr�@pTX�PY�GT��Z��`�n>ܢ	�����&Cc>A��X۽�_#F�=��
,+��U��>��8#�3�vv��X��Wx�!c�mF=��sD�_+����F
a����	j�^�]��FFaT(QGBe�]3T�ʠC�dNg�B\7���M�s�*�LHu�y�;�e�t�����C�Z�(���9�8q��O���������Kr��:�:	u:C�l�c��mӣC����8
��v�s�$�-(�s�h�����d������ϳ�#��J�殉n�|����S���*|�����*�ࡼ3�]ͮ�rC�EY�P?H2�pu��a�����Js`�c�:�4N��K�Đm�2�[*7f���J�n�����t"+�M�Qb|��ư��)e�ϰ�-`��Mއ��"��^i>"c�1UN#�;^�tZб7d}��/w��h�q�����[fDM�B�0m&C (�mWY_$,��a$xA�ly�m�5xX��t}0|�rY���^m�������⪘��Az��s��h��77?�^��z�i�=�l=���\A
��Z-�|= m�3
���?�I�c�����IC�Ͱ�-4����E���5�Q]�]��R���R�����>T�g���2]����(?G (ֱO��<1��wr_����u�ܚ�����^X�2ʔ�789� ���ɿ�U<(�?13��9���Z�D�5���A;{d\�K��	mÂ��+6��#����s���v�]�-i3��k�V�zH)I�yg����K$w%�w�Z��o�_x~*fg���o��6���u>��v��S�a��y�o�6+�:������~v"9��zG�G��J/[�޹b&��3	S��x�zvjؽ(�2��m)�2�R� kT1Y���c?���ْJg�-�$��^DO��oH%"��꧙�yݲٮJL���}�r言���[ۋ�����[�z6ڛa`hy�)���ɑ9>�h��KE���\��tgi<��d��U�Q(�'���}��*��k�2_ ��\���{=}=�E�`.�2Mi�5���Ct�nq�Gbb��KɋS���y���Y@#����g������Qg��{`�~�����~�\lډQe�$�w�ܣ�(��]ϿTC��>�=A*ܴ�ǹ��fמ�hO���iTb1����WAT?B���gt#1�p��`Q�[��V�B���G(����atW�Yf��aB�\뚪=�����;B���ʁX����B
xҎQ�+Ȼ�,+#1�������M���W��K�MP������p̛�8a7{�G}-��e��7�� �3ן;�R��_sn��iɤ}y_8�$h8��$��Ru��9K�sa�jP�[��*@��iB�*�H��<��
S�CP/tR�a�ń�?�Ө8!�ju��:.e���_��;&�b]i�i[�i�����h�y��z��(1W!P�C�F�n�8])��l�E���������/3�&�$A�	�1)Ɲ�y�VF����WA�I��,��L��يJD�毡!4��큙f�S��?�o�� 8�9��s?�Py�X=���)�8tw��f5d�VO�F�A�~��
Sl"�أ�bx���ys�g�s�o&T<���F���>�����}C������*�.}o���q\_E��u��
Pt��0�[��'����~̘���-g���]6�X���C7�@i@�︆���Y�g�҇��Z���b�G!��kn�����/�Iҥ�\�l�-EN����2ɲL�gy+w�Az���\�2)�gWXza�m��Xۗ�+��M��[2�A�0k�Cs�� C*�/����^E�Xo���n���{����s7\7�~>���Yq�^ ؇":��~�/t�]B}�Gg;7g�k���n5�HtR�����uO���H�\��Q�ٞ?���2�A��W��BW���[d_�Ud:m��A��b�B���&K���.8�t�v�{�b�d2N��O�}*�����	��$����k/���t��^�����I���2�w?ѩi��ZXO���.��*�wԷڂv������ܘ�KM�?M� ��' _y�[ma�+_rTG�)I��?ޯ>������>�el��ͺ�9�P1�K&�J����`\)F/ "j�,ϸ���]�ھ/���W#\NQ��YeJ�P*(.%zn5{VG���<se٫/�+@1��`vf��ᑤ���):���A���s�W28���\q)�_��lڬ���{�����?P]��$~������Z�C���F���53���H=�2|�殴�qa�<�̐D�>ôoNa��V_(��o<6�R�رtwy�g�^����51��J��6l�T�\a�5g�����K�ћ����%j6�A����]�S�;���[�a�r=�e�yk�;Gx������)�/�@<���BT�F=JV޴9)�q�ꂣj�.C���465�N�~��{�}Py��&W%�ԁt�Fi��w5��Ao�*�59�����:ə{�,���Ő���P�K ��U�y��[>�3���39 S���kJ�ڷU��Y�Z����8N��o�����`Iػ�R���Üz���+�B'(^_G�Eo�Q(!��c)'+�8���7x�R��G��JF��<�ps��y�4���]]6��0��Ñ��)��1
�5�?$�g�Z�轭ء�3s����`U���10�W�B��D�O�1�@��H�u��;�R�1�tu���%f��:ҁ:��-^�#lQ�������Ic/�6�e��!���h���uv2+�N�ۋ�ad%�w���y�n��,���{AG������3�3I�/���n�I��Q����)p z籊���_�0ر��ٝ��"�%�vr�ꠚ� C?�^0���U3�)��x˰Fɏ�M#}y��#p��Z(rf���ݑ}#���<{���S�8�yw��u��x
�m�q4���ƛ-n����RՀ2���M�=F�S�lgmVCT���ߛ�9@]�����յ9�7�{˲����f�l���������¡�ퟅݎ�U�'(�w7t�S̠v��������+����*?��h�½;��o�&���=�� ��_ a='��Z�]��2�g�5<<=��p:��(�p
K��_�0�,��헱;�^��k��Y��� je!</�6�%�G����iك�N����{\����A}�����(a���Ə���φ�Q�T��1�ӆk+��Ae�f=�7n(߽��&p����'�x�������7��T����@�H�gkKvmu�ضhj6vIA?k�����_��FVmI�bt#�� GE�vy������6u�(+Ai���FO%���:��F�����#���-�+5�(+A닉o�
w�ID�~���w͊��^�L�K*�g��^����\p��ȶ,{"��^���X��8y�烂k)��й��� _׹z�Wf�3ul����'m�;{x���r+~�ܲ,������d���w�%7��^���G��+����{����/��6����N��h̨�[X�zu�ɑ��D��9>��\�x�Sv~��XV��z���Kdj���u*�IN�0d�3�j��U��|D����V����_��Y��Q򌢴a^�CX����TU6\����A��x��!�̆o@�����~��כ~%^[�o�"__o9k�D`*v�៺2����p u7��́nf�f[U*���D�&�]Zz�{ʪ���HR�j'����F�R�8kD��X���?4y�^QM�W��AE�WZ�)�9�p��R����[����z_ZeS�qE{�ŷN�J}�T^!`��(o�l>u�`ԋoGA�3X�,`�fg�4U5�!�)򒗄>Ӄۭ*|�cT(Ƕ>��@|ƞR�0�ާj?-�������>��W��f���ޮ'��"��nli@U��l8o�S
��"T���n���w(��kҰ�e%$._2X0^��ŗ��/�pIw˩K{@�rWp��30z>�`��w���9�[�������h߯1���ǭ`����2�Ɣ�ڐlS�򶭁ٟQ&V�]��G���n�3r%��tyE�8.��U��� ��yUϺ%���Q�+�⻹��U�� ����7�o�G	Y:��$�b<%7�7/�s ���Є��,%�&�s���)��%9�u�#O��o�ӎ/5�
L�w������{v'_@���*\�J]���6���p�|�4ۅP!"��wn`��=,k��z&ܷ�S�գ=����t���Ģ.��f!�E{�������-U�7�,��+���[X9\bZ��_{󗸝�%Ȧ�.Cc/�:�Y<�o��|	��R|	�z��Lo(?�﫟-L�Q��Q����N~V�x���"^��גr������ʣ{���e�r}3K������*��^�nO�;E��X�3�!#�&�h��̇%o_�	�!0�����X�K\�뺆�	���(K�FY⟣��ˬ�	~� ��N� s?��d]�,��U���jL*g8�1���t�z����<$��u6w�P-+�,�K��\�1V�G{
%�����U���w� �c�º[J����]�Oo�/8�����Cp���l��Ycl�~&�`s�!��xV�}g�/���s#��IC�ߝ�I�B�{x�B���uE��LV'��f��4��j� =���@��承��p�[��ط�溤H�����/�#���-k�I�[q�?!��gۮ��㈮�4��� ����1��{$�-��L	Z{��Tǎ�tH
t�u�E��x������w�0ؾ7�~p��ا�^��N�r+�g�?���$�kQ�\m��{����Q�����k�e
������Ҡ�:�kw�S��-��_i���Y�LĦ����7���e$�ύ���<��ب����J�Xr�WÎ������M��b�래睜����!�ԗ1Ihr���|ex�&�'+Aqf���!wɑTvnu�#�$�j�pg�02U�i�z(��X綩d��<�?���Hk`�U~�cU�uvjx<��0���c��s<�G!�e��S(�?N� ��>�v�fe6y������� /ГR�x��z�$b6�WI��g\�Dſ�h��5�c�g&E+tx��w���,o�Jj3�!1�5�����W�,~d^��-�1�V{��j����뇵3Կ�bY�V���=���̼�>�-�Լ-��R�!.��9�R%KǹNO�-��禼�;�y�Ч�;ū��#�u���}s_�$}�Bg�qj��~m�J�%��J������}�������9�����,��Բ�S�e����h���tq� �
u��.ժwZ�c^�~O�ҁ�G|��[�����õ:��6�;�e�K7
�
�f�?	(��!�l�B�b�����o���ޑ���p���؄ٯUT��Չf�H_)�{����f�,R�Qu�v3训�?յP�>���G��_,��������U�NA�����k<9k>���2����� ��K�˿K��d��:V�P^xX8��87���ء͖{��+����uzsW�����D��q��e�{둕��!�pJ1�d���9i�п4��c.����.q��\�����|ol���A�BgZ4�W�(W�g��XI�\=��@�T)�8���N�'�Й�[�W�w6S��܁�L��ЛЏ�J��s��'�G8��
��)ª�$�5�W.�N��<��sJ1��.�N�J܉�io�B���[�S��i�ſk�S�yq���;���q�+z��ii��~$�������v=;#h��Y��y+ �6}u�ɲ��C�3d�����A�n�����N=-ۭW2���u���f������=���s4��)��_���g��~�-q[��g��v�f|_�\�����JP� ��5���$��M�u�R�r��3?�qGG�y-=�H�0L0�?�p�(z%7| ��N����ܴ<M@>UDB��m�sQ{���'E~��3i��8���=t7A^ʨ8���
�qYm�p9c/�B����ۆX�(��L�8��8�ڷ_�)fĤ�/l�5s�y@�wH��B��$J])�ԛ)�X囵���'i�� �L&��33�K92�I��q���=��fT+���bc��O���W�w��%�4R�%-nW��n����軌����3+��k\n���uj|鸭�wrBi�_ެh�"w���.�oE&���s�]�!��=s6q��A���D�zCAK��`�2 ~s-�Ι9�5�P��)��Q�r�r�N^���� ����~��.��H�Z_2�@���7�4��L
��.y��{8�\3��57�!�3�ϗ���zHg[nn�$�Z/�6ԔG��k�G~^�|�;�l��7�3�� %�؋�-K��|um�v��
���e=����q��Dx��	$k~�����/���ʲ��*BL�����
�
vE�-(>�����|Y��i(��_@:��xv�$���"�C�����Wn�榊�����:s�e�̃�H�e7��^m��$ʿ;���Z����m_'1�@?b����#}8�������X��1���H���F�Ia�+,Sy��^��T��CC��w�o�/�E���-p"8Y�-��@����n|����0�a�w\k�WF��8yVH��m�� Ct^-j	�^Zd>����H<��<��m��WxL^��Q��3?�1"�_��1�_�56.�쉮s���	�@^��"X�*�K�f���N\)Ζ���y�)$NcS����c�	q����H�?n�Ϧo��|V�3X��p�m�]�n�d��́�����*ob���j�?�9U�)������0|cxO�f\t��&��Txq�����T�H�q���8�#>~�m��_)�G̽�����Fp��i�a֩�φY�s(����Ƿ:J	A��9�7A7Ӕ��R�����W`��3	F�@�RqZ�)a�k�:,?�����R*��|��N
1����R�����%��� ��{I�Y���1�[��Z��5]�c�c��kBj��7!�o������Υ���5�v���Oi��Y�� �D]N5<ZA�ʲ	@�R�Exʎ3�I:L˓�9Φ�l���ײ�~��.U����-��CG-<����}��qRһG=ݬE0�J�ν~��H�viI?�ֺ�;!�Ȩ*�
ߌ����(	��{��U���3/�O�0_dx� ��)���H"�!��y��/��VRF��S�Ђ}�����̏�wLwhD���V�H`Q�nsQ��g\�e��a�19l�UD���8� �s ɋ_������>�������_A��4�a�4�yî}�zm|���8}�����+Å�4a�>43���m�ɒ*���u��A���ϥh��.�{�6�	�>/u|N�:PN��0'@�7`�v>C��W���5�s��A�/#�Xm����"��(��gA{;|�kŜ��DeU�P3y���ء��0)�Q�Lt��������վ�4��8L}n�t��;$0#a��4ɨ�>3����>6��'u�'�U_ѣ�P+ŽlY7��s�F9X�y���Hj�]�u�`���ho��yJ�y�1�!�?�Qub4�35�u��($�sL{�"(���2-��&��|��1�u���z��"P�H/�0�� ���/��
ƣZ{���ӯJ��c�[�����IE)tA��D�ߊ\r���*���3�-�TnI����f��.�m�w��n66�����`�=o���yy���շk���S@�œ��_-ގk����W2�N��ҫ�ʘ�q��4�jݘ��S��YV���_$#Ӻ�<���7Jm��N��ʽ���	�ΘbC��M��®�t�<��\�	�+3��S��pl�[!1�0�J�d/��{�&?7(�>j���KߺZ��~��u��8�廇�,����\�������>,
��-����e�v��A�yM{����@��n��6.��8��읔�p�~��*^х5��}z��w��I�PO�vI|�K���2[��6�JN�jDq�����s>��^���"�{����)���57�
�J�>�4��a�Z/�A�pC��?{i��qԾeZ��tm��o��p��|�YLw��a=t#zp�	��\Z�A�-�8�� G=��wc�=&Y\���B/����g�6���*[+�B^�G��RmM�"Z��B�I 7�}�4~�#��>DR.�x�����t" ��`�0%�M�	#'�#��S��{m�M�k{M��mא L��j���K D~��A߲�P}������|>�y^f��_Ȅ����:������_,�
���2w��ʥ�8���F�Ӧ�$�72����
�q+��� s�����=��z�qN��Z��?7p���{d��+�9寍��	8��e��|�=�_uo&km�+qC�
�����H��}د���.iD4,��GZ=���}Sv�Y�mJ����c��)MSJ{�F���	k���ő0�О��o����n�{�V�����z�D�Ck����w�]cqЯ�nȸ"J�2͗4����f^��W���!�ow����M�L��r�E�A���nC�R-���Q���5���Ehl���웲��p8�/�X̞up	��
��DO_�fj��Ɇ�V`w����^�i���B��
�I:�i��|�9܈�nк5zT�G����V�Z�YbV�YT��~�������
ň��o�NWhmWj��z.WF}F�?vx�:q�[��S�t��U�.�@�9�tu|8w�6��� �����Y��QU�+WL5����S[;rj|�i8j#I�K.��%�&�zD��Q8	�[�>�<�K�H��a�2�˃�i�������p΀�t+pe"�c�DC���0=O���	� ��Vо��5���X?��ƪ���6.�d*�6:-�#�&fT���b(Uu��+�s+K����o��hس�nj@���c�K�D&蒬��K�v◕F�`��<U�Ul�)�������}�_Qkw ��3�X�֯�$���kH;�-G�T]���qw������	wx��0<�Nڭ�u��q-[�4�D�
�M���f�wv@�"T����3=!O��т�wid{x�¼��r����y��D[��Mj��6��>�/��0��t\�}��l�B��5a�c$O2��ގ�A4�k���]$�P[������ܯ�y�Y�-4v���<qg��,�g��D�4�=$����,
�}0ݯV��jޝ9��	ZOV#��Ӫ^�0;e=M^��jCk�)۠<>�������>xm�^���v�ab��Zϧ�*J(M-���<*
�^����Z���&pO�/Y'F�f�h�
	���(�ӯ�`�^��UMCg������]��(�6��s��߶��6��{�fU7�o��Õ^���z���@�����nf�`����Ik�E��n�*_��P� ]ŗ+%�dְƇ>O��u�����$���GE�ή� �غ��)�J�i�ܤ,�V�10�]�F�4����-�ѹ��+WM��-i ��H�ش��c�HD3��e�U��0>�0z��1۞����y��hq��S*��˧0#`��3����w��t��2����H�X
�z�<ӧ"�A\���\�����C�8����������vv|��r2<�>�X>D���
/"�q��X	��/�~7b��	�֫�a��ղ���N�����y˵��aF�u-u�z�"&z�Q�B��`����M���F;x��P�	%,���S>���p��JE�>W�}�t��X�T���ɿ	,Ê��Q�}ءj��L"U[�s�e3��Q�o7ܹ'cK��͋_���.�e*)�_��yB@2I� Q�P��<O�)���7#�bw�p���\F�<��3+�g�GR�,,�<�[
e7�薆,��xu�ŭ��y��U阖�>�@۝粉f�����g�˟���Lh
�u�=0�O:h~��Ω�Y��;�R�eK|�*�h�lm�kA�у�����,�&�?���|Y���/2��&k�Q$U%��93Hi
����Nl[Lgܴ�^�)�� �&f�����$�YfrE��M|�!��(�LK�p�t�F�)�JG=���M�'�M���U���p+��V�qݼ9��ç�Q�~�3
��Us��6�t��o������*f�� ��Ӡ;�ڡ����n Ng}�0�H��Zyz����Hw��E=?l�T����Sl,^#�+4��I�����$���y�c)\%L0�k�a͵a�d$�4bIiq�jЖs�0h�������r�u��}3�*�ګp[��8i�a���F�2uRU�m@���&�8��Ec���(��n�j9�E"s��N��q�d�:�-��lx���ψ{�L8�~|�lCمnǸ7+��0ّ�y3�I�}�T����ދ+��?����?����(��Z�"t��vt�+�m\t��#y�����?lR�o�@C`�ݮ:bv�� ��Pd'��~������1���	�yk����r�/̂vɜ��Z>$��lt�u��1c�!�t��eVU��#�t+<��ECXbc����h|%��	l��ô/ ��?�|��-�<u%��u1<�����wc`��[�*�ps�4���SzK"9�E>r�K�Qb���\k���
�㘰w��`.���sY�hֳhi��VM�.���Eq1*<���ƨ�I3>���w� Jv<���u�z�߅}��$55���%�Q�I���	
P�f�w3�����g�l�ߙq͊~J�{5��71p���ZR��4�Jdb<,�0ۦ��r�!t����Sf�� 	����-���;fK�Y�7���n��9Pf5�p~��U��Qowtߏ�����h�ߨ�ƧR+U0���h1I͙3qq�E�=�׫%�A�ּҲ�fS�#�(�~�f�<��h�V\�8�F^�b�:�r�P��f�$N:�y򷞵e6z˦�<C�f�D�h�Yt4�%��`;��&3���Ο܏)�����"m�|�3:�r�w559e
6�Jճb�i����9<�\�����v�j~Fh:?\]d,�.��#Z���ּJ�r�c?�`�¶���ƍn[�����`���G&��	sg%�������V:����s3fuЂ��"��q�F6eBCi�і5̈=�>$E��ne0�]4*�$��t��Z�T�c��yܱ-����J/^&u=�p=��p����!��e�,����Hm��+c�58�J�寤�bA���!J�9�Ѩ�\�M!�Z[���'���>�@b�cu��sZ'��{� H�~���۽�<��V9uR�ɲp���чHJNS�#d�N�b&�p�T�P��l�\��!��\�F�n��8t0lڻ�$i^����]^卌����C���3�2CcMA1������xI_�?2O9']
p?������p5��V|4�W�ݝ�1�n�Iw�:���}9L�����
�-t� ��~�ͅ���ͬ�0+)�ܴb�}9�sV�;��۬O4��&$X�F[ƛ�T��.��1y������Af?��N+"�I��~S�Q6N�M����F��]��R� WKğ�Yi�҈/\n�P�=�D㚊��En<ڭkfL�nE>t � ����3�Ϩ�w�,kY�V�?��̙�.���Gy�p�M�u�t�7JH�!�#���g���'�%����y�ױ��ԫ���>q1̇�B �Abu$�+S'�{�L�N��W	���Z���]��LqC��y�x���*�vw]`�m
u���3�G0�
�$�~���W��}�y�g.�����2ieJ�g[�;�B5k�dk?�������^~����4�Gm�R��p���:e�J�L�+�y����z�ʟ���9'��xA��=�͇g�� T��ڽ&�(B�hàF׀t^-�o(�Q7{M�3!����tw�`׀b>~�����B0�9Кw��i׶��P�掀HzP1?�-��ea�W筮u3M���)�׃�A:�W�g���<^~Jq��I�%�q%�]�� �~TN�F�*�T���vso�E��:�=�@�1U}�EO��N��gR�E�	��&R������Z�ax5��$&ihb����{�	��SCUs���?�ǽy��W��f�u�oh��g�xG f��@����TAc���YpL�GD,�ڮ�B�J ��W�2�+�#���=L�ιY	㪔^S�?�A�x���6xp�M�����
����YoKL戇�-�o`�97i��4��x4�	O��߹Z����v&M��"k -�#�CӨ{KR70o,�)�����es_�N�x"ǼN�/5��֕aXTb���ZN��
���qr��o�d�9���y�e���'d��1v=�]"*�A^R,�~h�Ra麗�!��(޽i���G������k<v�@�Q�t*�uu�L����#����̟/�v�Z��a�pp�8��S��C� �*�c{�����
z�U���u��Qa��]� ��� �v�n	W�1��9 ��h��4RZ�G�9_�9�_ɱG~�IH�.%n�)��qb`j���޻kZF4���<��t��,<��F�$��:8hz&ϚV���N��GvaGlA�m��$���9����̒ݲA��}�fE�����Ē���CS�=�P8w�%o�X �i����/I�Z8���z7T�H�u�	u/U����U&��b$]>��l���Ks�/���K���1�_bmhy�<-O��>2f�����i������A���eʯ�⡢Z�TRx�2��������V��M/$��vCPe���:d�2bO�vu$���z~�<q�W~]�:6���9�&��ӳ��=�22�)�>�ao'=��}W�%���:5�����t��.����^n�z�J�cM�Ug>��5��.<7�n��MW�p�@OP~�+�*ީ6>0���x}�R����/��X��Ya!$p'ҰŊ��ЮI��\�Q���
�K%2.��=-4]p��h�ZyRM������ｖ�A��<�#�ppYc�=�I�S�	�֮Pq1�W9�k�v����U�`v��!L۪҃��4e� �C֖=�15���k��#\��R��dP gt�w�N������͆�Ǘ's�;���e��3`<�jl*@��xd2��Pa�6l���6�>w7����;ƨK�o�R�fp�5��^�%U�̟'q����Ȃ^�����b/(+j�)n=4��V�e���(�����9�Zzz ���:.�#"ݜ����u�̿���U�.K�!��
N�D�������WD$�
d݀��V�>e_�Т˦%a�f�p�a����9���'��y�]fKLn?��|������"8V���|O����T�7CN�U��ݑY��4�.�y&}COM,|MJ��ּ���tG��R=d��D�nʰ�/k����=@�f����M���"��ϰ=nW���_�Y"����W�!h����ݳ���2O��v�ԛ\>Ԩ�kJ��1�����b��egr���w�Ŝ~�f��+i���u�c��5)o��H��U��Ž�$���P�-8�[����+V:OW�]!�/ĻZj)$�_�W����#dH-%�m_
p#/˧����Z�<��T]�\tc&���E �*� ��p���$v�'7Z?|���e�[�n\<� G��T��7Z5%3�Ft+�i%O�?7�[2��;�%�����5�ݻ�ء��K����
��g�*��j�ۖ������Al�%'����BA�ڮ�n��G��1�����_i�+2�nŸ�@s�����I����o�'����J�*�)�o�=&���)�H����Dy�[�.��z�r�v8Li�`QC�FZ-N�2
V��:��mЪ��B���uY�
�NN���HM�D+�]=��ſ��	g�>�|���]/�fѽHW���CevҲҷ~�I5Y5�ý�.�& ZEi�[q�ev�wR����WG�h��b"33���{�t��
��i
������M>��/�Xqfl�\VI~��lm唸���,N�bg��v�,��f��-m�;`A���d��k�9پ7�م�V��Q9P��d\]�9��]���K>=��W��V�ꖷ�Dɠ��1��rB񺠾�U��[>���P�_������<�#	��Y���,�y�;�B��bψ\����c�R��Y��R�Je�LW3�y�1⢭I+�����Ւ97+��)jjE����jo�c1�%�e��gN���޷*=��w�@�'�T�d��Mb(暴�N�}��>��k�]�r�ԋ@~&xD�G�N%O9es.�M�.�ie��Q�jj��nc�0bo5�k�{��V�hgԮg6�{w�FD���WQ69�x��U5����+��T���/���a���30��^^`A$:��aʃ�8��%�����a ��ڗV}�8�-_H��s8�j��!q7�6�"8�-).��ܭ4�q�w��;lH�`�w�Re��������o�!6P��%V [�����-Z\���v�bg�p�+܌&;����xH��A�%�G�E�ŢS;�*��]N�&I^߭	N$�5b�F�>�@�����w�������~������%'��ܐ~�!�徚G�W�soŔ$�G����g#�%2�]�%�Q��D��[����n<�ޘk����
�r�
)��ؑ�jw�y�T�m�|�J��G�J�_ǋ�z� 1u����(��C�mY�t������A����2�䗒_��?�����P��k�֓�i�����eg QC��\gB>,��/�Bi2�~��#�Z����߃��;� �����1+��|�E�!���l��[y�t�Ή���&����U'E\",2�k��)5h�0�]���1��S�K��Z��Bk�z�F�T�y!C��&7���k^@�l�5w�.T�m�Ò��t<qj����_�'�=T%���@�uå"��N��Du##�6p�q�{6Ӕ]�Aف�]V����~P��1g�0!Lk���4�󀒣���:v����YV����q���d��")8�/ ^�w}��U"T�T�$�w��T��[�5r��B _��sQΤMz�:�Z����S�K�P쯇��3K��ۅ����K6��l�fkGA�?lZ�b�r�v s�]2�߁ϔ�����U��c0 /q%�cDu�����`�J��*��"-�������]wG��<�{�� �>�n�ާ&{#������{k�G�Wz��S����U�SS·Z�.���i�:HQ���L^
V�R������7���{j�ΈF=2�Dᙎ#.�Qd��;t�]Yh�p)������=�"_��
`���:����wW]��A%[�bO�^n�"	l4�s�\ٳ�^te{���z~x����"9#I��Y"<��	��jZ�)ů�B\��L�l� ��y���^Ƿ�1&���_b�;���)�^>��(��\D=»M����	6���q�@��c��)�����/�Ctk�b��#b��i����'���'���s�b�d3Y��K��@��37<��������%v�9��xO��{�Y�_3�k7GT!�ǀ��;��kj�J�1�r�G�_/��qy~x���DkL�X$�ù*c�,*����q�����C��yr��/=h��z55��6��%'C�/��)��Y�K��0�ܼU,��P��ʙ�� Q��V!e�ba}1�h-�w�����r��#"�R;/x�����]	�\{9d?BϚwM�0��2���[-�0牨�a��\}����m�0����T^9��}��+�t�꺶=��7y��N�s��e+� T&�د�駸B|�}��I��s����{��ꢠ�ּ�(>�˂�QS���TYh2s�g�nݿHg�#o��l�C�Kr۷Uxc���S<^xj�LT3�T)��*{��y�DZW���/&�mT���N����p��ڞ��>�Ľ3��hȂQ�(3!��c�|�!ǜ��	�1�|����m��,��Ϙ��zL�t�-��ɚ��"+�*D�c�����3�(N�d(�����v�����T3�\=���k5����O������Ԏ���}�F����t���w�*owTݧ�N�jϷ�R�?3k!�T�C�mb)v1�/�Ű�}�zZ�����S��oт�����b�-���C�� �m��>J��O��Hr}��R�R7�,����)8*����F;TMc�B�BUb�TkiA,���Ѷ�7��|�;W(�T�|ܲ5QI����B�����l��4��G~��W,Nq�0�$Ta��Q��%����T����m�+3��G�q�z�>�$$���(���F��A�%ڐz�I������<�5_��ִo=r�޶��,��?���V��_�0���l�h~+�F�Խu����wN6QOk�<��<qN����ep���åMf��*GI�6+-�u��"�k�D�{�$�\����=�ygC��Z�^�����d���<�1������w!��9ݪ� �3��;��ʽ��<� �-�O�?7w�Y:�o���?%�_�<M��S�Q�6�dT��Eo蒮�5WD�\C���455*x&��ZĚ_t��H�x�:,)��,�r{��z��h���oΊng~�Q����*﷪X��T�GP4��Yk�\b����Sʪ�a�7�����t�6��rϛ[�mJԺ��4�)��"723!O�����ˮ��=Z�E��|q�*�������������V��I�cH�嵽x~;!g��#��{7���M��#���R���ǖ�l�nb�� Ή���݅��.X��8f*a`*��
�wC�� ������aI�JK1�{,~��W;�wq:W��w�L���'�k�'oB�ӑO>3�3M!����M隇m�a�Y�l�ݤϋ�58��O�77���U��?Y�9t?3»�8F��
2զ��h�?��F�{�?��(���ޚD�l[j�L�ÉٗO�>�dm~<x�vk�[l�"�+(�"CwG�t<�X�Nh>,L:X���v�C�%�浪ϋ��\�������N_ ��ٜ35�����j�/p�^h�m��{d(�I�L!���L?+P;�Ny�;����RB�(��~{b�3���a�x|�����o�s�ܮE���r��)?���rI��Ka)G�ւEC�5�vZN�������#G&��g�n2n��{e2�g�<k���n�Xxκ�I\��A*8��W)-�"���Ec��*��ؿ�UuѪ�Dm.Zl���Y0�W�S[�"�dq/YS�r�4���J�/{��#QW�w[����@U���Q~?����j�9�}�'�3!�r#�eء������m�ҽ�X+׳��e�m?��Af�SfW���G�c�j�g�qH
��_��Jl�3�Ü{�k�k�R�(P_Ff� �5nټ?�VL��+|!�}"��jbO����]������o�W�u��Y��c��o�
1U���H=�/���}Q�w�zԓXv7��=%�d�Z��k\s&�l�=��vô=�Q���Jq@���;��K���y�/.����J.�'��~n�οiW��<%e���f�X�>�T�(Z~?��L�Cֳ7P��xҳ�x9v��W5��x�8_�#�W����p��Ibk������~ďęb.�dT�v�k�S�Lm�z��f��@`_��l��e�����jTL����;b�rt��cuxke���o�{���c����V��`��~���$ϷU!	��d��q�jdGJه=.@JJz6vܡy�����[-������}���w;;�ب@����WZ"3t�2�]	_�k�	�q���Au�u������(ʤ�ۡU�N���ve������gfS��T����;�4�'ǂ4���^�����r�?Ƹ���4`��c�%{$���EY-:�����9�SS��2鼝����(C�6Ky���>�^��'�u*lRb��$'�ePe|[,r�L���(+*q�X���2�.�Z"��p���T,&�J~;^���H�*�|5�Ǧ�2>Őn�Cͻ�C�HW��R8���԰�y�g*���>���FJ�M��Hjac�(�]f�V�K�dٖ|Gm@h�~��ge��GC�0k�m�PV��u9�rQ<��JA���@�[f�B��'TaN�p'�uԳ�,_��"yE��0�	�x��y:�C��������LWDZ�?I�:,��S�����]�����k+)��:��$����L��儶�82Gfx�A�[OzT{�|Y'a��M",�<�[Sfz� �ij0:��ͫ;H�sAV�G�H�p�!&���J-�z<��M�����xn`bpKqe7���k�ZR?��g����K_{(�������:ɾYM����Թ�v�D�5n��]a��u_�C���ez��g����#���(h������+93Q�q�Π�I�{ʐ5���G���o��p���2n5����O���P���pqC�z��h����~9��t29T�-��a�]��+{���a�����F�_��Ϭ}^�@��'}}�;��Q5�n{eeY��x��2.������E�*Q�}&n��Ģp�����u�<�_���#��w�R��'���n�\���^�N7]��D<�����������g���A��Y����_�W��2Ng����^[�i�<���/t�E��`|3��U����Ծ~e���=�������Ji�M]tJ�Sիq�č?[��\2��?�S���0�F�d���-��j�B�!��Bē����Ja%u���0x$��0����EB����w��K��'_{x�j�<N>ξz<��nW!�ٻLt$w6��)�h���y�#�(^i� SsCJ�EcE��|iJ��Y��9�S��݉��[~�_K����ez��%F�C�\v׿~XB��ڂ�?n��rI�C��[]-{!
W���5A8�,�gN�$��� �S��	�#���JZ��B=:`{�d�f%�(�ʬNac�j[�S�-��M����-�����Ű��ѫl3=��i����KŪ7�.!.������y��}�~6��&�n�ϱ �V%�X�{�����du��#��>�����7���?NG@���/��SK�"�2Cϓt`��޵�u'�C��F��sth�g�p�%>���2S/x{9��o�H�BI��1����h�vW�n5sx���E:��⹺�F�]��G�����ȸ��Kk�V��"���&[�S{DHm�PG�!�#^�bǑo�3詳�
���V�<�~$G�ߖl�o�w=������B���) ����|�m����L?�Kg�M��p��!����N�1���}�����FM�L�X�L�*a5ȇj�C���ԕ����4
�<U	䌂h-�Zo��.�xJ�{�����E�1��k�3��$�r����>��V*pOK��?� ��,�>dg%M�����pO�:�!�\�ӻ�$g3�,B�vӗ����ͺ�4�wV�G}%��[����08����&��zS�-��%
߹"�g-���p5�V�f�$J�~�hc��Ƽ���[�8����oK]�Bpi8��e_��־�?/�	2w>1?��%\$U������㋕����Y��y�]���T/qr�PD{�^�K��#�0�K��$�il(}lZ�v��þ�=3t�?��2���vj:��F�ǽ�D2ޭV�PP@o��6�	]iy�����!�xL,��E�Ae�? O���c��Ik���:��)�	K�hg	�8��e��oM�7�_RP�cp�����OK��D��5���m�W�B��KAU�~�L�K���Sm�&V���%K���]�'����4�u!`���s�Ç�7��0�Ŭ_�k�8o��d�����s�%���Fr+��K2j��
�*=�RD�qLkͬ�.���8e��U�b�%�G��{�;�O9l��EN�9�i�O��*Tc��4W� �V�}�Uތ�2�T���cp)!�(�W�ֆ�m��k-�����}��0Wt'
�#���_��bJ���~���KO�nr����qE!�~���3��e�ɟT�����I?5��8��{�;ߤ�]��s�ed�b��4�r�RZ{�fa��)���N�ZJ��^���ڏ��L�AG��	�x��+~ �y�;�5q�����
�-���m^�qG�7l_%OB�V	C�L�GQe����5VZu���jȑ�U��_��>��'\�al��^�h��<�2��,*3�u%~���N/��U�Gu�͎���˰rDK�>��c-�y�˻�FE�
��p���������L���,K�ݬ�O[%�3i P�ɀ�+�?��2.:Q���T���A\��$�_���-�V��o�p q��%[�|��ԛ�����B��sF[= �X�8S̤��ñ���E����ߝ�4~ᅝ��&�O+��i��ݜc�<��c-�Zh�/�aW^l'��F�nT|���Z􋿩F߾�wP��;%���N��� W&B�Q��A
�dd3�v��Ab�:�6�X>ޓ�$T"�(ì����B0������+�}�\=�%2����N��|��Q�SbкK&vR�s:K�w9�O��c��C����%�$���*등U��ٸAzI�̟����r�D�#_��À�`�aQi37���������al�e�'����>��� �T�ব���l.���3唝�>k����M���ﭭs]�X�w�6m��F���/��f�$M���=�2�&#*T��!�>���)l
Ye�?Gn+��!w��u?{r�luC��uٹ����f�4�譬��f����`�0q*^R��z���M}�lݾk�����m�:j��q|=��)va�&�]ԃ-W�����0v�y3�B�Tw�<�fb�t�M��`WCLZ �~(B�ޖsU���έ�a@s#+��ڢ#m�&2�H�zK#=����~厘2����L����YYK�@Q��:�uuؓ{%?�����Z����/�YJ<���R��n���u#8��'Sf7{�5�\ʵe�~xc�'z���y<x���B�'�m�p�:?]�ws�V�����n�\v����^�k�����l׬�'�?*fi'^�G�xP9�I�Tp�5�"L�G�o�t�s8w�m;��5��1fUy��bu��$��$�~��P�C�|��\`�e���B�g��K`g_��@Cb��c���x�׆��Y��W������.��J�.W-|�njPrL��H:t�2!u�A��#������[�6)�wm���O7�Z�z���ˋ�s؄����PK�@�M]�<,����u�p�z�p�V�>@��B*;'�����ǃ�i-���OEfj�EYF�x�[<�p�Vn-ss/D�L�(	@+Ty9 _K�*�|l��ِē�}�hF$�̥���v�z^��j(�(��qc�r���uU	a�y����o�����JDӆ"n�^���#e�z�Š+����OT>��U����GIu��`H(�Z^=��ВH�,8 $}D���á[w�����4�Z�&&��w&T�aַO�.L��y�#������i���X�sd�~�9<�[g����2mQ��yP+��5Th��߀��s���ӻS)�r��En������
��q��OH�(<��Ow��m���	��H�uSJ�~ݨ8��2OAd�$�/�Z#ok0�n�\g�8|o�����7=����u�M�	`�}ӹZ+%y[��Hlwu�`�,��"�.�&���[����?�ܵ8XWOY��L<W7e
���{8���M)�Y�
���}�XÏ�o�z�0�(�3�ڟ��ѳ��J���oh���~��z�����������}9��z�T�{'|�dPj�0U3�MB?C�6X���l5�H�zrP���] B��6�L�=Q�h�pF�/��b���p7�&8�H�-,��Vu�������4��֫����|�šM�?L�GBE����0�p����K�����P�DT���إcZ��R4���[��F���eTi*���d�5"�:S4����S|S�!�և�[�?�2wy�)ōJ���=δ�Tg��V��g}<۾��յ���SPD�����#��L�z1��m��v�a�|UP�g3ZpOړ(��;{�C�[̪r�â'O���pY��ZtFFG=�?��A@��q�I �.�xX��~ֿ��o�%��44;�*a�>�w ��N#m৿�B��]hk����O_�8�ktB���|ٔs��,�����Z� ^�� m�D��Kho/X����^P�"q��L�L^��;PO��n��tG���7�y-C�-�7W�
ݨ�	r���m�6U�H~a\���ݯ�ه���w#o�Xe�cN��ޥ���<i7�Ӹ�q��t����̣�I_Ğ�{��^�����ˊƖ�.�|C]M�ޓC�	��F�����z��ҡ'�F���UQ�7����ޕ�R��Qj/&WD�9Z��`|�=Ҧ�o�O�h��B��UZ.>x_��}��}�a�y�
Ӈ�<a����O�Lb��%oǐԈ�2��0\
�B�r�g��K�9X��<��l��`Vw�{��`��تm$�E�+%��b��T����T�c��	Y��*؟#��ْ�?ޗz5
��ϛηu��lߵ���p���S�R��h����~��� �5� �΁�O�]����CY�m��x��8�C�8��f��\.��"tJ���g�A�\��F���z�$=�4ie�~�MNN�+jD,��f�s�,�����Ĳ��bj��^ޝQ_$?³ k���IS�N���DE�x��.�6
T^RtuOQ%*Z%G��\�+��Pq�i�"G���d��.^��[^�˖+XQD�uJ7�Gb��lFV���t&���nxi+��۹����0KR��a��J����~��7�m�*d�ѥ��G�~�	��W0B�XoN=��iS���Wn�x�����{�Զzc�d�gI�՝��U����FP O,��һ���F<�c��J|�_"8(���YY����I�`����]�"�1R
Ҧ�P�@�k���<n��S�M�:�fyc�hT�ͪ��y4^+[��,y�ȯ3XgzH8�3Uf+p�z�kR�2L��I�|��M@ȟ,O�gĺ�����Ĉ���j�;��=,eF������XB��rb�h��Ƒ��s�a���ý2�޼���e���t�k���s=i���9T��� M3�n�\Y�^�]d��l ߍ��B�srθag��h.0�n��lwV�_���%�r�vuK���z�`r�����s�ME'�����Z"k��ʂ����Dݖ.�+t8)btiR�C�턗�hUXi�~�3=�j���o=���F!j�����ۇ�u����P��_y� E��H7��f��z�9��-�2�I�:�Fw!�`�3v� �_q#�`?�/��f��X��V�Das�3u�d��J�'M�Z���DJ�����z� s��En��z��1�}���pQ���C@������-f�
�4�}bϿ�X�VYM%������P��7�b�����w�-���i֫��Ul~Cح���kPL0<\��p�'���V�XA��3'q��k$���밚��S�%����������m-�6�~�C����C׺z�+VF�6:����q2TN�y�o˚u���>���u�"���E(�(�;��m�M�-�l-N�욇�;Q�ݶ���N��8חp��P��3��Q�A�ߴ`����݉�ղ�i'�y�]����>�l�T���D�2�VUʊ�:�?+A8������_����l��ʥ��oJ���a��'8O�J6��pwN� �dŃ(��˸�\�������
�Zq�z�.s4��ab42Tփa���c�.�9h�ٝ,�I\'	��^=a�2���~�"-N�P=ӗww�}�[#d��*x�ɅZhSVl6cS�U��*q��(�� ��� ���g�/
�DAG�#�w6IϷ���
c~�{fv�ߏ\"!�=!U{�W��v���jQE}��V�(�#� ؠ�8�l�q�����R\/�.1`Zbt(��D2��[��3O����/�|�e���i�*�����d�ӏ���A*��W���f�>J�Ӣ�	�_n�퐳7@O!3�]eD=� I����#��'q��efQ-�ט���J2�I[F�Ν�����u�c#k��<}|��kx�c&@���;� (�nZq��#����^��Ѻ{�v���=A��ΪX�4z��]��̮�{��Ɋ꫒�S+}�F�t�Fkbϼ�E׈(�t�@*�Z�����>�Q:�[���^���y"~��cJ����=��S_����ݮ$*		�B�˾�l#kBd���-{�${e��d��"{vc����1v�S�������s�u��:�=������X�C��C�U�@�Ild���� �t�D�R��S��Q�\�τЌ�Sl4x��N}���9U������_ڹ%R�!��~�a ��?�믬#�6'�oL��
*!�=��w~���k~ZS&zc�!Y뜗������a�&?$��G�ͭE���a�,���
A5�"�Ж˵~w�h����׬gx0}�J������ݭ)+?o�TA)�q��U��}p����A�4F�������`�=R]�te�4��R�]r䴁��y峥���U$5E95�n1f�[e�El�?֫���д)g}�͖�}g�'b�W`��K�З�b!��43JR5H�۱��
��q5�8t�TC�+q8�`�eQY�[�:&)�9P2]�X��<t 5w��ƿ�s/��f��)��;�5�n�h��t @���mȩ]�Ɲ6
�m��i�>y|�(rJ���u�I�d\:v�r���Yv�x�vYG���«�
��] ^?�Y�u����]F��v_>�(z5�Y��ݲ�-N�y�fh௛����,��e���\k�@�!{@ۓ� ��u��I������]���a7�VE��@�"��Id٧	�s��Va���K�bz H���mߥѨ�?��Y6�{z�;���0[s��� 6Z��Z���21�y��B���iV�e"� Ǩo��������]�Ыs�bu"�ܿ
J�^�� �04g���7v_k�#m�̦��k��ig1(Ԉ��i��NI.n��d�/f]�ܟ� 9g�eCt>�x��!墿��kX��m��&AE�9T�BW�D��HF)����f�x�{�hzNo�k{ a��0o�Z�(ʵͳ��a�8q)�l^�J�3-���[�,AkLf�s�o����Ķ��v�B�i�qg?�����$%*ϑ���%��HF����t��	)��Eco�b��.�K%E�c�|d7#����l;N������\\@�_���惽|?;��f�����0�R��-�|g����\fnxxʠ�2��pJY��1��ƙ�H��P��w�++@��%1���uS~����Z3Ɩ0D_ӓZEy̡�x�޾��(�}4̋�3M%�%#�6�왷6��ҘS�
/� ��,���� ��!�D���U8=W0eNDz
��~��ZG�b���/�р	k�Ը���W���'/_�Ř�y � ��:��*S����d4�+!���,{6�/�:x�-����<R�����Ա{:�p@�3U�c_���/r��O�D�q����#��F��;��x8���q-V?�j�"Y�.l!{7�B׍(.�,O|����ǎ���i55g�J�Ƒi��-
Y`B�+9���#��T{�8��� ��/�^�p�- ܞ<\)u,/�;ݙ�L5����??�y�<�Pɻ�|IC���B4����&WZ�D@_���Hٓ2�B2L-�h������N�u]ij
��)&{y��4���Z?/��y��t*ʸ3�yܗ�k5���v����� 4�h��3��o_d�QgL��n�ݰ2HZ��B{fn���Z5�VE�Hq��3 m��
O��mЗ�W��)Fu�5�����`�� .�/z�Ӂ��Ys譺*F��v6��H���g$"f����RI����(K�OΌݨu�]�����j�
��;��\����F�	�k���J� t��kP�u��ñ�Y);�@�'��J�G���Mo�v�z�~3��-׵g�}9���)��3],��ވ���@F*~C�ʏ���2n��9�n@;z�� ��A6+�۳'j�X�\�&�:x�Zpc!��FOP B�x1Z�ؔ�%S�"�7���wb�ˁ�$��ߏ����/�\����[�{�.�\�,f#�K.���w��B`3�����	s�����W�*�E`�ޜeϪɆK�f�F{�B��/H�w�&�<�n�o�<Y�9�~tT9	�5�)=b|���ߠ��w�H�Id���e}-����|���0[qΕ�֡���t ��J���$ꏕ]U�?��	�Ʉc��)y�ys�T��eo�B� �{�'c��:��Em��^
�M��S�-v��a���v�ǝׂ�}��n�aа���=<���I��npf�Ǒ?t[(���6�Q@��9�XC��-�R3�����g�r;����Vv~��"^�wcfm�S�X?)Nf�]r6�ҞLk��l���hbto:/eYZ�9�r`��זP%WXX�#Ɩ�F'Nh��ٝ��G{�A�j�c��_�͟�&��w�Vo�C���a}���N������"�#�ձgSvZr>À���U]ʽ�ï;�fǗJd��8#��'�ƿ����Ӹc'��8*���a�(����k]0iJD��@F�w˷�ձ݁O��+3�c{P���U0�4��J�B�R�j��A��.��p���E�}5 �Ž-�K�΁���;��&͔��Ə;2]���E%������a	{p"��r�	��-[c�o�o�ىI;e�ٕX�խE�l�>'�����Yr#�fA1�UU���pZ~�3 ��.��-�	��m T����g�P)�݀��i�1�_I-)T*����(�ߐ�f�wj}���	)�0�G��hC��/�C�����vt���C6�F5<�PĞ��?v��3�y;�⼕<
��R���g2̒�<Bn��H�=�X/�2{��TK�98ٔe��W
NN-G9^����ϟ�ZV;���(e-�~��J�+�t0�t�ӛ�Pr��n`&�Yc.�ҽ���QE�3���ˏ2;b�W�1`���&��<?��tx�y70)հ������N�,����lb̻ZK���ՠ\,:�9	9��pPD�i�c3��2��jM��##����ٰ����U�C�n|�ErWS�ٶ�����j���4�+:y R���'��lCK",��\?���mg�'l��3a�ЬXhK��q�5��f4��I�m�����p��7"OzW�Oy��>�-%�uc�{�E�t%ҏU�k�I�=	�sŝ�?>HT{�
�o��\��2���F��[YZ�Y�N�8S�7o���`�~|���8ǸNV?�oXz�WK�� ?�R_Hp��Ċ��3�JԂ+�Q��ڻ��}�������#�9t�X7���<��W7fn8|�3p��f>(t���
��9��?M�O�����6ۡ�FO�$�-w�C��(~5叹r����C�Բ��ٖ��0��V�!c�5Ln9�ь�&~��E�K���9�KP��Wϫ�±�03�:\գ���8l�R*UpUG�0s<��|
��v%�D�;���!D�R���[&���E?h�[\��?�yS��˭�Be��1�n��A���H٫F�4�����a���y�[���%���9����"	S�X���I�)�J��S��K�)��_��g����?u�9,�Qb�s�ǒ�%�*k�x�D��6�ٸ�����z���~2�����w� �9d.mS-�"���{b�Vu�����34a����&,ǂ)Ѐ���?�k57��?	�]1Xs<t�q�rϊݟ���/��x�6��h�;���Mm��(��>+;���r��KNN3C9�)��'�*�
lF�I�!�>����Q2qeUV��#V��+`�F�_���
���]��3w�(��|��������sNנ���l]��{d��i�BI�+w!E<:%=l��h+ROy ��\W�B�2��#��"�m��q����=#y0yEp,2ܽ�+�b�'~�.{&3�w�N�3��D���Ū����,ͣ�r�y�
'<�"����?�$�_b:�_s�q||?�C�+�yGg0�{r�.�_G��Ơk����~E���}��S^��L��i���ɾ_�\}U����p��n,�o�+^x/����ahJ�b3���F��"`������8�q�
���9��xi�PD'J��q�P$�<���FMC����"���S,��)s��Qr&���H�yx8'p�C�\"��g j\���<RH*�������!J/*���4�e���dk�ϙ;+R��H~5Ho��������:ʯ��f'�"cu$͊�w����L�G�n����#�y�5.:�>�@��:�ur94mo�W98#�'hx�M�v��v����N.,�'�7g���,�8�m$��=ợ��^ U�eO�H���z��h?��XG��2ㅘX�01���߻ocC(/�A^�X�\X��=#�?�w���(u�>{�Q̬?fٳ���A�?���>���Q7m�p)�x�!%��G
��B�SZ:������W���������4��Yg��ϫ6��ƛF׈^�p��
[ :��EG�J��\Ad�U8�~��m�ChA��-=�]�@��=zzҒ4C��̕t�M2��0����" ����_:g�,x���3�����9;�i�޳��Sˊ��;� ���q�P�q�g]b�������k��	�L�!vCp��Q���c Y�ghז�i�D8Io��V��ܴF�����j#�g̳>���q'����:9��A㟽�\f$`�>��I���NI���'l�pe<1Eh�^�[�o�x�.����침Z�!ĕbc�S湀�G�=���
臡�1����6Ww�{\�v��>���ʂ�=a�CI_W�ʽi}@�m�l�9��e�ު��W/��~Vu������t�(�.�5n�pj��[w.�}(8�u	�gɓ�r�������TZ�x�)>&H~pc��fV����`/�}Yw�k�w�r����u0�ޡ��\A0��f�.�]��/���6yS����-E�^{I�FƬoO���Ԡ��K=��hT,�~&�ץ��U߅,�+�a�m���a�z�+�eݩ��L<���s�+���j(�HZ�C�@H�Dޜ����oq������C���W�F��� �ާ��V�%][q�Y�"f��;�&F�Qy�ָn?,��� ���E6Й�6uK��)��?��-��aS����!G�D"s�����g;f!5�v�Q/�J���[���M�Y���ȻZ����J��&3R7}�B�	08�>�;m(�o0�I2�!}�{VB����|��LS�@_Űӯ�U��f#`�Ͼ���>�D��{�S��ȃ��}�,Š:�y�q�$��(����I����4���_�Ԋ�$�fӍG��_t])��*h���w�G'�z����� �)��A�R�#�g�	��naiل2t[ܪ�_Zq8�g+�_U���Ea�K�g{Tm����[g�W�;]������Yӯ���ͅ�������3T��R����T��K� BL?�$�V�K�G���FP/7�MFא�#���c��bU���?\�|��H��1_l�'��������lxg0�lӟ��l�2��+Kq,�D�X��w�u1���-Ǿ\�)���������X�5�]�AW~È��ݍ�R?]p��7�S��Zi���,UդD��NX����{"�\�t\pv-6�μ�>��n�����`6K���D��^i�9�F�y_����=j��k���_��m�������7Z/)̨�M>	�C��K��M�0A]m�<b�2|B4�!����ex]Mzn�>>c]���ah�5�0 �t��Gأ �Pa���P�3J =�%�����_-�׵Yy�W�A X+���!ho�T�Npʌ�㝰!�vL �o�+�ĥ�1P��f��� 9Y��ƹ��ȅC�O%�a|7�"�Z��Q��]D���桅��~E�tb;���|�9.k�̿�ч�ņ���~_D=��d}���a[M�L�0�z6����t���̭�������o	�p�sm����7���K��g�&MC�Kt��!+T��	jJc��T3%n~,��k�^��g!ؔ�s�T�;h�Q5w��ÿs���[sս�˾��/��Rz<��2���\�8{�nL�>��_d�U�y}t�GC�B!��k��̭�J�K�}��a�IoʦY�_��=� �������ͫ�2�U����V8
W�N���%p~>m��A���~��?#�^|7�+J�wJ��U��mBU���u.甄Q��h)3�v8ݽ����מ�UM
���}�N�䦔C�Ҝ0?�n	V�	��S�����~��Y�Тf�"�=c��S��V���a$�)��R�gc��|��w����C�k)Y�#γJW_S&�k%Y^�
)1���B��*� ����f
}��r�r���F֚�z�<,�d���oؗ�D�zV3���L��&���k��v���HBYiU�_w�(�aWt~����ҽ����ڋ	���+�FJ2�^	r3:K8f�4{BPջ��[9&���i3l%�Q���?��/���C�2;C<=�Ș�4pD�(��=�����tgW�#�����W-W�t[C�Ĭ���K�}G��F�[��>̢T��K��EĊ��2��AE����g�e�2Ӄ7^4~�_��F%�o��r�/(�q���hU��E�%ǭ� ��Gz�5��O����@�f�'���⥙"Lȯ�
b�qЂ���Sd#>�:d�B'�&�M^"h�=x�5�7�v��9C�D�L�å¦�Z��c��V��m(���|����Ao����^�|�\��(M���s�ǆ�,�����#\�{k��<�IQ��$��q��QQ��9F�}k�N@?�V������댢��Į��|IP��^��IO�u�&Iϐ����z�Vr��B� $�����W���M�^[$��vB�{1\g�?g��9�dp\��q
�3K�Dx%�%2������:4h�^����"9':"̄���k���M�Q�q�Oemv�"�&e�2p����l���We�5t�'(s��~��y�-��H�z��M��,�!'m���u��2ơ�n�R��J3���ԥ+��ʃv>�7+���n�;;LE�\*��ʮ�O����6�Rj~ї���ݗDf�܍�Q�&�4��^p�r�i�æW��'�w�7?>_*J�"O{�1�6��%�� 9AhF>W�QAv;O5�yQ}��ж\��/.gVʕ���"�������}��`$�\W�N[z�K�4Z�L���qHy�#�7A���{��ߎŬ�?Ԟ䉌o���NT�*��Yr��]C��$�ҏ�0NH�S=�#y�~>!��/���3(�Я2q�y0��p
ݶ��pw��^}�����Q0�s%�{	V>j��o���[E9o�Ы:��
��a��� /��4�������]Ik�s7�$����z����CG?Ƀ����v�V,�|X���5no7���D�a�im�ͪZ�����o|�wQ�!Y��dB��Y��~,'��#9���!���O9�#��㖽�$>�^��vП�x��h�8�$�VD���&j�y�������Ҟ[�|��٘Ģ:�Q�Ǖ��f�*������q�v�S��"��m%2�
M�b,%*�9�x�,_�� �G�����܄�xE%�3�Z=��N0��:�vCz��ts��jA0bm_�y.�u�Y]�\���7]����A�����CX��X�J����Џȉ4m��_Q��{iu�ye�;�'�~�v���{�K9�{?y��1?�/�t~S�:4�ƴ�d��q#A�����t�-
gsv/�Y���,�-{�DW��=M��YV ��:W�*䦻g����oP�q��M~��3t��-{�����طA����&����Ԭ�����?w{��]��s��Ikq��-,�o��\�Dw�Ԍ�E|��H���c��~�[�@�G�綢(�T?s�A@(�0�wgX����Aߖ�=��&u{y�2>N��{���ڮx�ǃ=�AV��lE���Zx��!_ӫ�}~�@�٥�N�W��	4�<7��5��d���4«�uo�0�-w�G`e}:��&��]�QM�C��y���㰙y��0�1ɑ�ɽ�ݩ��"�L'�?^�Hg���G����3`�&S���m�ؤ��L>��~U��_Z �n]	:\�i�s�|�HZ&'���[wQ�~^�޼Y��i��������ߎ��؆��VǾ��s<�a���w;I9tm�k�@�siRN��ۻ
�U<Y9����Bp���*���*�y���q��0��z{'��z�����E�T�����H(�Ƿ�u��}��~Z�F�`s�Nٳ/��U��=*�,�Ӓ�҄��~<��WL�G�.X"���l}W�>Ǩ%s�!�7��f���iP�k�?��x��������.[@i��z��6���H�]���<��,�x�y�����u��k��@l�E�&���q�oZ��c�uSW��X�+�Qg�`����\��3�L����j�vS<��7��>0�d��1�y�v>�,�<���v֘�^���;1q~\I����,5z��+t��K��
V�ۙL��XB�s��I�]�4��I}Y�r?���_������%�2�y��?Q�Od�=�v�K��)[�濵���I��g5�֐.X��4)�[(y㻭T(��=(}�%���Ÿ"㯏�ܩ;7�r/���)�V�2��	"�ju�}f`G^/�|��+c{�G:�,��`��G&�_�[QWǯ��}��;:�
s�{�J�S��3��s��Zm�J��mQ��%'�_VX�;���@��'��)��eF��ї<vy��tK��Q+9�xq�E��j#��]9ރ2\�J��뵛]8'�wL� ��F?ux95נue�Ǽ���e����f��/��lX���(g����@�f�J|�(K��q]ۤ���qe��3ZE�����ݰ��]����^\�Z4lW�8�赏�Uf��o���0e���j��E�ޠ��m@Ő�%�ǀ�Ti�:7���_�c��A��!�f�˩ιoSV�K#��{[��UMk�L���"������Ǚ�_����SP߾�Ln���Ȑ�7]���"�Y���s�������\y�f�f�g�]|�����������'�^�N򎷕���-|F)�i6��Zy�����'�^�q__q�T��(�����>�=� L(�^�O���j�(m˕gJ@+��
aӓ)�)q��^4���z�i5�L,����=���AA�$��b�u�#��e+�G�2h⢆���P�I��aW̺��a<�͙3����_E�q���7��Gy'2F%n����?�>��e>���r�N�6�	�E6���TC��
��ۡL����z�ۥ@�\	���?/�д%�-��8�3�o)Q�sB�:��KWFؤ�t�UL v~��H�A�?\�0�+��%W��>�;���Nh��[�`O�Q����..t��9x���]��
^|/Z�K�1�c;?��̙�5{�-�{f)<�V��Fw�t���f�O�e���WW~�\G�D杭���tT��|��v{��1v�3����2<��PØK�	V�!�z9�,�����t��7L:큾���g�K�� �� 4Ӷ�v�.���_r$�b�r���|>�)4�ݕ��;�Zv7���-=������F�vhUĻ��-�Q��>�f
3���TT�%g&��/��R�V�[Km2����%�v��&�l�a}_��n0�H��c�!�y��]M��.�`۴"%h�T��H���a��׵Kqo���A��Ӑe��7r�)������0׽�&�m������m��I��l+�����Փ�LSY�� �<�9�{�h�����y$n��z
�TOv��ݶ;�N�J׺�D�Q4:�U��x5�������P�%���o�vz���q���@����zl��!M�/g>��d��v�BAI�c*@s�����/��E�EBS��#eD�#c�K8����6�w�����*����i��?��������,��7Gԕ�O(%��~:���kx)KS��맼�:6��!�1 N%���ZS�#%P��EY��t��Ƕ0�aOP�kq�͹-r��\>�����5��]TRo̻-->f���~����x�}�U� �L�}�΅W�9� �i��7V:ٓ�Z�8;~�3�������N�@��fNTP���:���AȄ��fI��,�D�i/z�F
u�=b�N���TJ��)���޽���C+�C ��˵���~����3
��#�ߢ���}_f�v��w|A��m�E��7� ~6����o'��L��0i}K羪Îe3 jr(����+�|����N"�1
�F���N�����{~����Y������&F:��r��{�H�=�,&�l4�D�Ɓ!uE9;Lx6I��u��΅��w独?[ցe���
�nǶ��g>��%�;���c�����"**� ��#=��y���AT�sY���-ᕗ4+���z��J4!ԧ9!�u�j
���nwا��Z�U�����_l���'��إ9S�񷲔�R��sρ*e�s��b�k��wтb�k힖�q�kjr�9�4�}�E�E������(7�O��x�?��?Sd���P�4��Цx웴?&�{{�x��c��B(�a�	+<�Jc����.���g�k��
2����ڞ��9�nd]��~*�j�5:���vz-��~m��2�N
����\X���1��k����b���Zmy�ٴ��UX��R�k��iRݍc��JW��Hߡ�9�cK,���o�������r��倯�_�ViY�>Ú��Ѹ�3�;���I�"�/��[KYi�X��4��[��7�*�װ��vh�b}����`��A�2���u���y�����ՑY���;o���_{_5T%]��a��"����Ջ��|��
�	N�W߫	��� 'Xd}?W��r�4����s�� ov�d:�{�Yej�J5?3��cMp�Jݎ��t��B�$�N����b���J�Ӛ��?��2��tR�/kϪD:�����p�).���4՟k(taSһ��)R�ODe�-���9�������}��0M�D�d��؆��i�ah�ff�gGŧ��n���{W	ފ��~j�ެ1�x9��RM�>\���M�z(F'�}X«Xi��E�%P=�?&>SlYw� H�I�j[x��Ȝ�̕ꦱo�q��9���65��QCB*�����T���]2�����i����zG�
��>�
��0�C�]Q�#�r��v!��d(F�w��X�uE�ue�S�j�~	wn�:���FO��epJ�E��q(�b��� ~���#�](V�̟0u����`�?���m����Ԕ��`Q��A>�M��3	�E���Yr#�n-B5̸���)pe|x��h��Ҥ(H��ht�|�;C��Ea����4�P���P��PЭ�洵��K���6T�Q�j��-���J'M's�w%����n�hJ���џ:���j��eu1y��)h�2��M�U�E>��4��B�z|����{��vG����N=;Ct����@͇k?8�I����x/,q��i�9<���L�	/���~��*���TvE�T����U>��2�P��2j�aM�4>"���
w�YÞ��!�M�Z��"��|��[me|�&�[᣻=��/�M��ݣkh8z-.Ӎћ��?��}l�f�}Y��x�}2�B�Y|�T��Y�W�g1�"�89�t�2<;�+�u�^�`��9�1"LP�V�*�gO�����I����𷞎{E�R����v�ˡe�k������s�mY^n`~�V$����bC����ͬ��6��dM��H��������������r��-6z>M#��Qr��F�Qd������J�g�Ҧ��s�K��^�Ұ��J�<s�h�^R�o$�,���ө����4�k��a�*�����[�b��~���b�˟g��*�`X������� 󏒂Ф�^�w�z&���c�Q�LG��$��{Ĵ�S��z@'hf	�[{4,�	C96��3MO��vQ�Bs� l쬿F�0w�lH`�4D�4�㏉F��Q%�G��ٳ$<6�Eq��ХtPmL�����r�V�Pd��N�.�¤'eVhx]�:�oVBC
�l�2�y�+&�g{o��tv_�jsv0֊N�B���$Hl�t��jē��U.rZP-iv٣'2V8f-$�+�����FQ�f�9��jDA�f$����T�w�<�*�X��9��9E~��J\O���J!�����/�2u�Q������Ӳ���}jD)�������|+�+����Y j@B��	���YT�ݸ��6��tI���hB]��s�#N�V�&S+�~��*�!af����q=Hk\R�Յ3�������'�љ�� �/ݮ��;�ׇ�����AK1�f�R�	Ǒ�WO�E
��7OE1�v��&<�{�^����6�'GN+�0��t�^����[~+Eփ��K��~��:�����D[y���j�d~�Q88���i�=6����;i{*�����A����Pm�N����U���IJ�6��*��+S�g�#)ώR���{�(�(�.�@��eڴ�3��hJ4���l��V��du��%|��薱��Db� �������C���_BOm�?�x\�v��"ᶓq��όM������E��u�����cX������[��M�8��l9Oo��Hi���T��D�)��	&�
p�h}E]�j��F���/bld�]̵T���;��%Xú���N��6���`vû6D�Z�ⶵ#�&r�/��V�D���	�5cSg�n�*����+J�J�wQ����q6В��{�]�ö���5]��fl�/�]J���5��p��i3��m���~iMk��s+��C�ƪW���\�>{�i�V{t�U+H���<
p'c�	N�}��0[�;���H��~�"6& �
����0��<e�< Fbu5w)����[w���
����uB�ic@��,�|�!��5��uJo��t�J�fUD�ܮ[�b�Z��MCB�٧�e[͕w_?��l��p�f9��pr�70gi�:�[�<\䏦��s[�	 s�}$�������{������J��^(����~��Z�R���o*}�V:S�H�7}��-�Y����>>���A@���y �r���~)�r�{L�IG����L����K�+9;��AT��CkWw#��f���\�]	]�J�n�c\���}6�{aȩ�`����!��;b�T����@I	�3LW&�ϰ,��w4��٩1����������i�s��e���a����|S3(��Y"��*�n+�틭-���N&��J�ŝ���s�����Jۺ�:�YnK:Y��;+k2Yx#V}�'J*n[��t(���:��^lK�cK���S�9ٮ�f��(�}Sw�
t��k���M��Y8�㧠n�5�������g��[Y�!�뱜���b;e;d�#h�_]�9�mm��4��c�QS�� ��ݕ�����)�r	��6uu�!o5M��ޘ+țӷl�-��"�8?c�3s�:�M�H���ﻣI��c�e��A����~I�����_�Vg�`����]�3뮴���f�r�
%�0;���Ub�{cz�R��3�L���P�\� .n�	e^��& ���������o�ۆ�س�c�y�@1�UY�����������n���Ŵrs2����_���'�����Q#�p������f�[)(�sͩE�S^��&�����Ҡ���l$�B
��/����s!��V_W ���������bk�M��:���6
g�.�`��#���8����n,��x�&�{��/�
  �����#6�m"�*e�"9�m��O�|o�l��P�^�)�k���D�$R���)r�[�I,-��'�מ2xw����j�A^�}N-�Qa�=P�0�t	�d��������g0F��c��c�*�5M|*?����5w!Ř���w��x��{Q�q��K�Na���}����k���V����}�𰬛�zU؜^7Ve����O�ͼ���%�C�$���{}���#��&�;+^y2�xtb"ywW9�v��O��O��!{����	��~ڬ�/���/�����m���9�Ic����Х{���S�=�����Te��V��V�λ:��C[:�b%f#`�7��a%��Z	����ѹ�D<Y�(Y�
��M���; 9w�7C|#�{�-R������[ڴ��0�b;�偬ρ�
eN�h8	M�g��OGj}X���j��L^Ϭ��rK�g,s�p���w$7m��v	���J�_u��coD	5���O�d>��Q�S汹�>;&���I����}͝��*b9sɀ�}��~��$��F��^Z�Z�lE��X�64��)!�%5����+Qڏ����O����~w�L��=0��k��Y�yD܀�;5��-���
��cJ�j3(��o��ɐ���wk�Ȃ|!1��l_g�ϧ����}�T�rgF�4��lVS/qcg���+���X7�J�υ��g�օ>~�-%i�Ҳ�kϾ��~%B��!�	�B�����F�JrQ�'��7ɸ������tB������i)'��}���X�=�L����j��V���: �Q�I�5�q�{�'��������*���X�+k��ɬ��y�)�T�# :݌�� _���I ��Yͦ���>�&:Gw����_�k���6J :rm�����,+zo�S��.h���!�ԛ��
ƚo0�bg�^i�)�� 5�k�0�S���5\������b�������rcQּ����1=i� ��m�����n����-)?�q�4��F��'AuJ/�!�f�|R���o�X��7�m��^�J8��~��7z�_�Q�0i��?���[G%��j��z�Z�r=���z)�f�s������4��q1"$�,�5	o�VEN1dO�����@4}�e|��~�q�4���x�,.�>��J�K~[co�P��b%~1����� _^�u44�?�=ǹ���_��0zb��go�a����/|���Z?�{Y� f�^Ċנ(���s��Eύ�O���E�=EZ󩏗�J�Y��!�	Q)�']e�8�N�!w�^X��i��u��:V�S�F�G��3O�c��C�vJT�����Ll��۝�े�5���j>r���Hw;y�+��/��8�-\��E�CWYi7�#`^��(�8�%��}��{�a�n�q�X�7�����'���ؓ����dU?�ӓ=��y1�.�j~�^��%xu�Çz|{�D[x�P���k��x�nNڶ��[)����1��P�z1���6B_w��!��[N����T<V�ќ���X�G��Ɗؚ6y$�c@�����wm��ɦ�O_����=�.F��N�y�g!�{�L��<!�O�[��)~vn"{�x�{��������'���Z�O/��F���^�1ђbW��1�I��غ�x}��d���~]8�q�ܩ��;�aiz��ZY���urr���-A�-X]���Ig�Oz>�J�e�8�q͛"���d,�!CZ��1��Y����|�S��Ϋ
���YV��~�^�pJ.ӿ��%�����)8�Y�Sa�[<�"y@�c�QC��7b��	�qW;q��i5�س�W��� ���u*P^N`��s�Fs�6�>#\w-v�Tڂ3���z�:!�}���f&<4�s�G�c',<=��f�v�~���J���Z��$�]�����s�����l,�zH��b^\fP��Z�q8l��x"ۖu�ɯ�oU(W�bf�:H�T,��e&c�n�uJ�ɢ�x��
܉�w�K�<�\�D,���Mdٲ�r�� C���� ��s?7ݚ�X,����]�*����
�c��;��;M���!j�u�����)Ǟ������ڶAI�qGp�Or�<4�����e�Q�R��v�e]���WG�=�����琑�o2����mٓ/\��A4��D-��y��w�.�UuuXt��K�Y_��ɇ;I��u|���?Yu�z�X4�i��n�PN-�^iw���!�c���,R�2���،��a+�%���c��^���1e��Ѷ�eGN<}��br��Z����\��;E�{�ъ$ӕG���"�S��E�-������G,����17ç`�NS0wi�W�429g51Qw���϶7�zRf�� ����0��v�P/�ލP��h�"^z�Izd%`�r'i5K��~p(�����PN�9���ޅǓ�m�*����阬�t�%] գhݘX���:�������󫊄 �ؽ��س߿5����D�:�4��Ze*��]���8�c�}]G^���J��x�B�uJP<��/4e�¦S�@!� �Y������G:�
�ou��3hE2�}cj��)j��sd�ֶ;�2YB�Bh��;)�l�qv���{(���VD���q%��oV"hh�!���[P7B����@��UP^[�G>�eJ-��11�#�!PKM^:�?�d��tT�!#`���/�r����7r����e��p�ɾ�� k]��Lj�XN����c�8�d>P��4�Ε��܋{���bc�}�J�u%������{?~<Q�?��$�sq�rs��>6�n�V�~9vJ�y��/MD�Yt���*��nz��R\�*JZ���L��9O����x�ء Ld:����	z$y.,�	\x	K�RB�$\lY�ɪ֊`�:j�L9>b�6�&I��� � fe��U YuV���"7a��܁YJ-�X��6����['kdc��q��_��CW:��7�q>)݂�3,a��m"`A5'QGg ��U����E+�=�^CD��%� B�FF�FM� Q� �D1�(�{�2�����{&����χ�����{��^k����&���̝����D�wJ�*��G=��ƚ�)%y�L����h�&��MKV�I0�acƻ�Ԧ��~P4H�Px�Iww+�(QViM��u�O�[�ަ���;����&�<�ehz�Z���}|�@���J������c
>�b8�Vl�&̜ɚ�5/����a���à���f9�ώ���7E���?�k�*�xF���X|�:J�����ן�*�~ndFt�o�u�<H�}��nNn��U�w��5*F9�=z��z���50W��lJJ�4���C۝�M�m������^�� )�M�~�����\�ۦ1�UZu���N
s4$CgC9�3��M�虼�ɔL�#�o#$�{.�kBwCĠJ��^d�z�h/`x�y��5&�3Z�Ƴ�g��^:�\�y�Si��81�t�����t�h��.�,ވ�dy~��/W���@�Bq�F��E�6��/2>�͏�k����L��ZQ�4���@u���D^-�M�;�M�VՑ9x4S��7���
��t��ϽX��;jRQ���~k�S@~��8����SqIVzc[z��S�p���D���I�wΫ���R2z�e"�N��w���U����9�	U<�u�?�j�չ?� �X�9�3��%�	"U/���E_tQ��,R�U�^�'K��nI�k�����s��7Mk�ctn����`�8%������*0���%G]��;�U?&;+��&H���^�(��!b�{:���)�#�h�G���a�D�(kn�{����<>:����g��`q�4X��� �i�}@��k�
]_�PRK�u2�����s���&�e�u{�)�V�'}�mQa���C�*�(��:��f4`T&�A�7����!���)�s}�)u������p�䵶�';���0Z�a
��tV-S�K@�k�;�_�d���%4�"��[sv,+-k���ԭ��8��W�r��ь��H��v�aޚ^��#�-=�D��§�)&�ˌ�f�I��WQ�I��ɚ��h�~X�Ov����N7%�o��������??�������E�*�Y�ﯦ!�z�V��^���P��cY�@7M�(���j6���H�@|��u��2ì'��\
��Ƶ�o�02��f�$�T��ƶ����}_�[Q�x���~���N�᳓�O�;����i�PT��UZdZ�΀I�|���(ngH�z`� �>�
�M@�%`\�T�Ս�>
�W{��2B����^��7ފ�i�n�ɚ}�}Hm���}�=c�Hm6z�)�>��@���V�!j���)媊�Ŏ%�J��S�V�P� �сTm������i�s�ɭDթ2	�^����IHME����³�%�dH��gD���y+��V��*�&W��kϛ��yT��9�~X�4P����6{��fL�7��t�m�%6�95�@y[�^
�:L��/�C�����#s:�S�HN@�����B��yƪ52(��xh�t��7����Ҧ�|������>�`�{q�4�gX�"*L�|��@�6e��_�aѣ�T�T��'��x�7!��q6�ǡGv]i�XO���K}�c�V�{W�A�%z��[���o�JK��.@����ʱl ��R��=mz.���`}�k�*�nS�W!=f1����7�cv�5�)	r�V��/��<5�M�9R!�9�h���h����5po����8N��#�bZ�o`.�Ǘ���}襱6g���Pj�ց�>���	���;����<����N{{���T&~(ʫ�ѯ,2C�lpF���49�����Q,�X��Q֎	ǩ�4��^�K�=��
�W�h�*p�ϛz�����|i�M#�n�.F0����i��������X�<ӧ�~g,���O�)ƍ�m�iz����H?Gf���ɲR��j�ö�ߢ�?��ϙQ9r�n���:n�Z�;ëN�v�m��}x������_�F�ΰ��E9�䢤�~�l�ʺ]�?�|��ޜ:�c���7������1[�TH�0�7}4w�3ǆm���H���/v�,�V��v
�?��@�5��l>���\
?/��C�q��ö91F���52��3si�m��xS�Ў/0�����L|�V�x��p=�[��-����u_I�J!��\}�<��20��7o��L�;(*���t����r����m�5��9��Tn�)�<��;���17�������Ֆ�N�(�D�
�,�t�;�Y�^T���/Ɗ^�K_ELw�t7��>�����-����>����P��b�/�o����������r�:�A���bҽI�ߡ�}C��d(4�� ��!⽯��zZM�1��)q�����Y�o��v���+9T��D
{������,MJ��t���9�P�Z�,�bU�q�44U�$@0屇�Ԡʂ߇ r���R�r�{	ɍm �W���g]A��F��@8�l�zolE]�z+��C覎�LR��v1땹��FϻLP��;ݧӛ����P��
c%��YE�=J�zK�˛n�g��yZ����*����V�z��n�<ڈ8R��p?P�85V��uɦ��wBo������[O��_�X�4�`_��Kr�:��Ɵ�1����ӭ�ow��P~���in�+cX~���v��\&�͆, MwX�Z���Zy>/��e	$M�����:��N�; 3��)V��A�?N��WGM�b����q1{��#���`x7�Ńtf�a@�:O��mh���^Y}��"U��RV��iL.�_��5�S��������-.*Ldk ��;�b_������Y^ߋ�1N��
��ʳ�� �����e��/������<�bkkk��o�E���\��g�~�?�D�*���F9���s�.ƭ̺,pAO]N�,"�IىC��s0!��p�+��X�2�Z�Q˲h8�3�
�����WII��^���j��D��
�D��\4ZR_<�RR�H$J��p�g5]�)���Yh񼟭%]��%��8rw���:�Y�2����o�)j'��o���<6U��ͫ"��/v� =�~�V/�{�&������^�l5�~b�ؾiȟ���M=�w2�v-Z��*?��$��W�'om��e.H�N�]Ww�J�,ڣ���<�^���#�7E|�mME;����"������/��°o'VW����y��nJ^��̶]�i���X����\� ��e�'�K5��g�=V�5���J����������c	%��Q�e%_Ѐ��[W�P꫚�OR+��F�2�ţ2�j��l����T���K\��E'��)I��Z����T-h���gu[n^=�c�U�G��祺\�����PR�s��E�ξklxPl��鷽j
"�f�>����w5��B;4���"�z��w�v�a���Gd,�\�f*��B�'J[ge����S�^����^=SG�$����������Hw�D��r�
^����*�B�����qz�=�'us30! �ς������v�Jb�N`@�Q9k�9k_pn,�G���~U?�]]eG0(BڥT�a�S*�|?���TI[�X��#��a[��^U*�o�WW]V�������Kb��8c�N_V�B��j\H�Bb4R��c;-zӎ���8��U�Ŝ�,$���O���'oqw�1��z�NI��EM������2�S�F�Ѩ��R�Ţ�ڒ[���s�a�pK��� c�a}f�@@�u��$px�P��Q[�Q�9û����zeff� Ī��1��_���Ω(
d|x�3L���2��O��4I�:q���5���N��6��ym@wOV߽u�	g�1+�C4�:N2#���p�۔�G�aA�C#Vi�F%�����
e3;�9lX����|��`W1rJfPw<� �L�Mbw�3d�:�8w��C1�~ҿ��_cO�\�+��9b@�a�͞�҉��Yв�/��ؖ��td�O��^ת�e��L�0	�I�	�
F��{��C�H�nG����][m'GyݹI����^���ru��}j��_��ѩm�c��w��v�w�^yd�K�f�j�w�sO�Ы����������w>v�\"e�|��7��m�&�����7C+��Ss��~
���� ���������)��$�g���6��GY_p��xr�������퍅���0�b�N����~����3B�K�Sr�D��h+�Y+ �(H�>8�
6I��0E����q��!�!�w�5�σ
W���~��Oд_��?i_�z8<9���!�%�ɏ�s���S��6%A�;ga�zQ���'��NT�ԉ�S�Z�B�E``a����1�Eer�="���7S=8�C�.��ǣ'�t�|��`/֘w�2�3Zi�p�F��"����D�֯.�}Q�X��ۇ���d��f�8�K��򆷐î6��]]Crc�͋���,�pw��K�_S����$�H�J1�qx��С�ņ��I[B��A)�<���#��Ы�Qq�jN�>e���3���Zh�/Bo�֏O.�+V7R��+W���kX���?�:�$��,�u3����Xų����GeS+i�/s�Zc;M[���{��pS�R��"���kSb���eb��|��$:�4o�ݗ���TwTƧn�2ݧ� �3��|�勋�R�,Gv�ܳNJ��5^�Qu����O���˒���ǟ��纎�b���,��%�L��xށR֤��[�iq}���+�U�F�L��Ǟ�z}��١Q��9��x���@�7�ᖋ���R�&��O���+�`���o���{Í�}MlIk7�eo���W���3=�>l��j�R����$���ࠛ.�ݣQ���$=�H��͖qw��$��ҝ�{v��̅O��WYWON��'ҭ(5Ik�;� _�޻ݮ���^��&�N�J94���(�*�֧2����A���g���K�|΋h����R�a�L@ٳF���[꘸�~��!m���e� ��@���_,�@N�g�Y�@ϻJa�	\�<E?\^��Ն��Sٓ��y�H>�{���Kl�g�ύs>�j�h�>4����b��q#L�����!��g}}^=om��G�^�����J���x!��Rx/N�x3薛��?�~�u�q+Κ��&<�p���^2�K�4��`�\��q���;oh����xh��~_��nߏQ�N6x�F]>���d���0TCc!k$1#L���4,n˺��(��7z�i�>�8��_0�x3����o���?ʹ��IՕ*�O
^�5��C^��S�=��Z�g�����,HU��p�%Ds#S��r�i��4e'$J�σ��M=s" ��N���]�����/��n54���Ywj������-~jY�b�G*��k����8&,��7t�Ѱ���U�07m�DH��`ǫW���x����O�c~(�)�)$��#�E=�<�����dny����*��t���W=&�n,��;���m�K��J��]��P�c�FSj��x�Nfq���q�<�PLcԫ.��:T�{���y�阂�}G�f��.ˣ:�uxrb��:�SK��.*����1]�!���Gl�/-�Ɉ����Է���4_=}�x���k��ׇ�������>~ ~ֳ�K�J��pw��|PS�t�7|[%z�%tU���_���Cj��1�۵�Q��*������V��x�"�~�H�^z�T	&b�-�qe�����ۛ�O��︃i8}�>m':lh�Z���Ѫ\��#�7{���_#?6~�i�Y5�|w���?OA�ߍ�ٝ�� �����z�v�Cy#�������d����G�D�hm1*�_'iy���fn%�
����~����RG�����������b��d[pYG�'��"D��̚P��l��r�à5�j�@m
b='�Mњq:�x2�������6N�/Y�d�8�eQL�3m��_J�h�����u�9��1�An�/�"z׆]�ܨdS�b�����+�Y�/'�Z���~�2�3�OFX�%_lÆv�B5j)n��`Q���9��*��C��*����ƹۻ��o��_}�T��w�u����Y =�g1�7&z�k�Y��LԶ�P_�T�\g�cHAګ�����CL����I&. 4�+�-l�	�C����;;]�s[��m�/;\�{LyMV[L�1�х��Ҹ�H@���7*��f���Ύ�^G�-F̠�O�l=��y�CهV<C/�����_@�_��d�M����`�J�F,-`������v���fT,w�k:v�]�z�Yn]}#;�U�A��V���*�罡�R4��`�[]U'����1wLf�y�,�~Sj�d��r�D�	Uv�;�틑�����Ǝ�	���cW�<����!��r;O�v���������ͅ�t_�9�D� ���x:%M`��"�� �鹺13+�LW���VE�I=�R�����tw���M]mގ\��>�g���uI�Pؙo`���.b�� @�F���.(I�C~H9#�����;ث6��k�y��,ZInIu;��F��{w��#O{4��e3�"~�'�6���.;���V���6����C���oGgp����8�v&�y�<sv.��d����h���7��Z�^H�I��i�0�����|�Y��SS��֭��%��D��0go�(�h�mp"n�)C�;��gq��9޲����c`ǵ�3��
��I�Rn����3}��>��>@?TY����a�
�z�v�ŝ�'�� ܲ�r��_�	DY��6A��%ϟ��׹2�3v��qj�}�6����������Y8x
5��D�>0B
	`�����Z��"{��胁B��9�P��󉚜�ҁ�k���MnD��<8���:f���8
.c��^��:߾1�BɡC�H�J{4�=urN������W���4^���:C��3�Ѹ�1音|��,"Me~���ᢛf�?<;�1�LJB�����78��]/�b�\-9���Ͻ=w11/r��ҏBx/[{�_>{�S+ô�=5��VB��=f�g��z�,��ܙ!0P�&���I�
�t�dE�yh� H7��3�WPĄ:�z<�qХY>�'u�I�v1�/. 3���{��r����d�f�%f����n!�Ĵ���y-v���ot�tD%=(^���Q�ݳ����@*K����o�����\(�QjY�Q��V~�t6c3^'��#$Ww�F���7�Mﶴ�Ӭ9Ffgc�Β��$qXD nh�����4v��� �o�b�캊�ץ��L?�)	���Kÿ�|.�߻�h�m}:z�p·�S����}�4C\�q(����w�U�5dV�<�F9kؒ/��il��~Ӈ3J>��m� �E5g?
�K Cw��5d�X%�������2	�����0E��|[-c��Z`�?���1�8�2����u�W�{j/2�[.���ʁIUė�F^�����*�!H�(J���ˮR�>��f���0KO�Ң��D��-��6��=�fKR�0�w�&ˬ�����;M���^sn���Nk���h#F6�o�w��k�rU�鶘F����e5{��Yѿ!�5����>L�Ԍ뵆�s��<J�@)��)���Fe8_�}������������~�f���O�d'�,������Ɲ ����˘�b�˝G?�)�y��_��t�J�nT�s����W�
5��J�7G�:��p\X%ޯʗ�|��v�ˌ\/��="#L@A��������I'B�[j�)�0�x���Mu��(�}fh�dH�����ճ�)���ȝc��b��嗗�2�@r�~�a� nM���8��0w���n����r��9�)GG3�0}��ɏ��.|Q��`Wa�Jm�( ���	7V���h�r���K?�0��侜2���j�HΝ�7��Ư`�h�j��P�0��9AZB���rR�K�䐷*�US�~���|O��/��pU���FT4�9Ŧ�P�BL���5�l�{����ҳ�p]�	��n�ʒ_��N(%j������l�;�?�_>���&��ͽ�nx8.{t���.A��q��m�HdրZ���,9{�yrʐ�"�ɨ��	�L�l�a��-SF	����p��!�㊪o$����7���a�E��NR��,��B~�����;D�> o;N�(�۔� ��k����]�n/�
CkX�.$�]x��U{�Q�_O�y��9���h��0X,�Z5Z������;��U�?����yG�*�,����d���gF�@�VVB���f�ym�g2|�<X"���[�#���D��R�]������&�z�O�z�:��`��Pw�׏�z�?�$�, �����kۓ�ma���0�3��k%�bF�E�(�er�gv[�$u�ۦAy]߫avO	a��m�]ZK�ky����7U�R�1�h�K�UTV��������k�#�C�Gq����5�� lA~��ks@)nsՕb3�p���8����������p�����5��Iw?��0٥#��@洅D�Z��c�����ӈ0�V9���΁�@�ߺZ�\D�=�������1P��MIz��{��'��9�x�tҩa?��ۥa��S�ž+�rʣ����H��S�Tr�f���qP^�3ɏ~qţr��C�\�l��(�3* Ҳ@�Q���t�LXj�;H譟��cc�q`�s��x3�U�m6_o����J>k���RD�Ĭ�|�[m�w�-b2���I�o�-�hg���>�yկ'�TB��%��W�lw[O1{,~��y��\!���� hbݪ�WPJL� ��K�ڀ3Vپ���R�/��6�M���p��<ڀ�g��<�C�����ն�Cnv�%��k& O�khqXY��� <�'{��˓�i��8٧즌2��߼�^�(Ơ����"�o�&���l������Z�\X�BCƸ��3��&VP�-�!���WoU���.3ɅXN�y�M%*ՠ�o<"Aޟ����,]!ȧMQOS5��ȳA5��8q����UUc �����;���e��j���d�	��7�")�Sb��?����֑Z�s?�=P�N�#�2��)5>�������aI���F�Ib�s��t�*Jr��n�!�P���^<���M
N�=����۟�6�4�RBL��Ef�y�Z�x/�o��L��3F*�:5_y�Y�t��A�.�	*�Z�Jo��\Γ�67�'�H;�u�w$@�M)���JP�D�������<Mat�?�_��0^#,�É0mGOC>�n�3�n�W�3��o� T��[Gmjſ�sUʇ�xks7�8/Ԧ�U�����I����������<'%���_�I届ij���}�t(��Փ�)}��e��f}jy33&��l�3����Gܐ _i~���b4Rt��F���Gc샼�[BR�v1���-�O��QcѨ�-��6�u�%x^��w��տʣM�U�����o%���N��;�����Q�ڹA	nzm31I˥�o���fJ�<��y�K{��#uu>�ɦ%_�_���N9wl#a I�Ҥ��H���d�5T0��@쉕��^߬���5����i���6�D��lu��I��hS��A��)� ,;^�~�{3�ЎO|P�ǆ���( 7t�N��� ����T�x�q���Gf���x�(_���%�J@���b�U3���� ���G��9L]!���E��Uo��-����s��J��_�Ï2��+�p/��;Y"���٦�j0%'���`s��xw)���,Q)��֛P��Z/�豯�̢���e�z�@Z/X�bߦb�]6E�t�c�M�j$�=��Xiܓ<�R�M�{�ak7�x����5���d�-����zO���(x��X�o��1�l��O�R`&ݕ|�*�z��+ȝ�]^��*@����{�̧�����e��5��~�H�q#I��a����*�\Ed�SP��f�p#�5*MH���J�h��4u�C*V��|�&�N���$��dd||��ӟx�������g��2;;`���V$jOn6��_�ƾ-X ��11S���[!-9G�\?�#�y����i�Ɣ�wP]!����'zo�]�����An�>d�ߍrT�~%�����`L�c��Ph7���06�I_P��f:h(���M����eP�΋�
895E���"�G�8E��H%�T��'��;>]�.� gv��l]喞�����>y�v�D����vV�#O�'XUՌ���^5a�h��1Q>o�3웯^��q] ��= o�˓�(��7�)(Fnhǂ5L�-��>��:\[������	������"��`GX��F�����C��VM���]�
VV9L�I?�M�u�b����i�����=I�1�ПJ2�d�͚gw�Ԟ��F.�-�x�qK�N��nE�O�К�.��~�o��vɋ<+��_R��rU�����E(tL�l앾~T�����C*�*d 8��Ch������O��]�Xf3��5��W2XO�����_F���.�nTC�|n^==`Ԩe&�#ii�wh���Bܬ�v��Yu߭���O��sN4�����h)�Â ��=�%{��!�O�x]��B�� ��mn����U�wH�!�5��ܔ��$�X�x���Q�fV�5�V0��W��
v0K�=�6?�ٜ-�q�(B��l�B����,�R���7:��v����T�H%Q(��R��0�	�|hk����tk��j�:�d�5M�b�~e9�,���8�8��]�%���4b�ޚ��3xA�;1�t��E�^����e�_ =VgRz6���� �Дi��I�r�w'�8�w���D�d��Rɀӗ��J}�Jp�8���J�=]�X���q]c�x%��uW`T�G�Jv�� �i���q���*fXkƵ������Ų0M}���uc���ٮ��t���*�Y��
/��5�z�������}.�m������)N����/�|:���I�aO��:"ט߮��|Yv\���W�Gw�z5��w�S���+Ot ��d��[u��\��@;Y��tx��Ʒ�sSl�\W�;�����|͖�2G|���B��PR�oo���zlll�9�yN3-j�9Kь'"dh�mh�3���HR��D��<֩�s7��6�#�S��͏��cM'��v?��S���^�AE%W>A,��
a�<�R���6�^��*Ӽ�eO��Y!w��L�x�׫�;ְ;wLк����{��t��8�&;����(�.c���|[`�w(ĽP����EE�HH.
���ny
���xQ'Hc���kf#[xoN���S�1�󱃈���C2ҭO���&�D����6W��3�u�|����_ً��D��m\4�Y�&_��FΜ�u��nb�~��e���DO��W��_�G��k�IzF�7�{I����JM����Z>��F{��C�U�5^�����?*.���hݡ�URR�eo	�-G�*, ;k3��Q��(���j�Q��S�ta�z����D@�m�����"=�b�ѓ�f��S%���\1��1�,�q�.�-����jH|���ꪄ� �j^�W�g[�u�x�Y48��
���[�l5Vj�����ފ}��-M���]�L1ٰ�擡O(��m�w|G�Ff_r�'���o{Y��6b�00Iʫ�NNF] ��#�G1�/ƂU=�,<��$�1
�:{F�n��fyQ����WDd�,��i��}6U��D��΢'Y�X�d�K�|��19V�֕o��VDщ�:=��%
e��9�8_knZ5k6&h*.&nI��H]y�8'���7 ���O����h��ŋ���O�}#|�6�A����ǀnY~t�E�/I{�K t�i@)��L8&������M�߶@���ޛ�9C�Y���x��#W�7�)��\�i�qj���-	��o��Y�7Mֶ6�q��ƲD������0ܡ��cO7�*��1	V˥�w�K��j��Z��0�ޔe,Z ���� {�^��6�FJ��I��ɜYl�
7����ok��)����p��>]��{��syTΓG�k8�^q����Yi���:7�d~��:�����ڟ��R�HI�o�wW�uo)���j+�r���*
� ���EJ�Z�4�+����>��y͖�y��mSB��{���>#
E-�[��8JH�x�U{���m �Can.v���	���)y�n5�);�����zY��Q�	�k+�[p����Ǔ���D@
�����Nem)5ad�LY��	7�*�.%�xa������e�ݠ��E��Ek�[�D���ԻSRN�pS����Ɍ,�qv�)h� �,O9W
��!�s��n����U��/m���m��	Y&m���Ť\0�?�z�'��"!N;8R�Y���s�!?X�[`39070L&]�G9�-H!j�=�n�S$~�n�^���Gg;m�WO�A�}P���z��d�W\p�/��m�Lc��umꌗ��<�!��fX�`�����
OM��(�Ռ��L���V�!�l��+����/�A�0�n�jzu�#�'�"3��<U�OB��U���*:D��ϛ2�c``@#��}U�9�=p����Q��:%=`clN�w�0Hn<�~ qBJ��"��kՎG%w����K�mE`a"��͐�㆛3�E�Ѥ�:���l����R��+{�3�I1��.���)ӑ<��P���Q7g�7_�x�q��[�re\*����c_7��
(���M���q_�B8ߐ�D�a�tĤ���v��f�E��n�KѤ8�m/����+��y�d�$��=��)�@��w~��b�l<�5ZW��v�\8�,�jy�� I�9w���7y�k�j�O-W<x}��;|�!��e%>Ɠ���:ш�,SWl��ݞ��S�ǚ��:5zx��_�

w�|���JWo`Y��p�5�E+@it�k��q#2���9X�U���S���+[�oZ�~� ��Ksp�3C#�-��-�N��]wf��X����R&b�M}0�5ވ�T���w.�\M�����8;�O>P��0Y�1�!�z��xi�B��U��[�{�QO�K�_F7��$L����%��2+��
����T�η���K���<��heԆw���΅����7��/�o�	Ҳu�Lh���ͭDW`O�#��%&P��Re��! ��%pp^0Ĉ3/A��]��p��M�{�!U7���O��1%���BggM��O��JDm?)^JUΨG�"�(�g�J\D���:��#ݦ'������>mt.��yZ��9R�uU�49|���lN�2�!T�������va,y93�r��;<���#�e�� ]�� �����S��lE*�:g
M�u�W�Vvz�jA˽:��(�r�Pm��a��jh"(%C3�m� ��v�ҝM��y���H���z�Ѹ�0����)�+��,Y冊�+?�yB��:z&�+L�؏�a��-+��!�������̑���ᱱw�;�C��<T��H:���۳o�Meu�*�OD=h^?ư��6���~�N4��?>���g���{�E���
�Zϔ�^-Y�|Asa;��K<��,M��8�z_W��Q�Ե]*Y�e2�o�R!��w�#6��ւ9�:�U'&��ŷ��Jؠ�4ژ߿��N}&,L�5����Z�H�y��FI�Bꣾ Co����[�i?.���$�����H�N][[�g�7S����%��
!��`���:�6��N� -�Ȋf�ObZ��8�kG�9VD=?�Wt{�+���9�q}-D�ҒZU��^ɔ_�
��b��U��f�o��ԛ���Hg�YV����ɾ�t���Q�zrOqYb	����^�96��7 �Ặ����K�eLMt�����K�9I^ܗ�W­���~0��Ճ��d#��1R|GG�ڋmXv17�iÚ���v�7�o�%E��������(�%�|V�-$���D�0����wEM3�����O�wtV��i�^�qGY�ɫ�:����:���T��5"Tf��ZVC��R�?r,I��3�qo�y5���۶�^ ޒ�%~I͡q�i�9�ף�ພu2�K/3"�c,�l����m{A�GQgL�R��# nBS�i|�=O��D"������rx!����s]e
r�F�a\
�Zۇ�뚶�H�*�3�y}K��Bf�R�(��s�-�X��Q��J����7f��n���'"���{
�K�ȫe[��`�`�z����P��C�Y�y�f��z_�u�c	��j:C�b-�|4�8V����'U"Zc��7�����0+�6Z�W;��;&;~Ԕ�{��Q���lb.���
\N��`�Ɋ�J�d���"���/z�|sŪ3�SS�yj�L�=�:n��b�����L��IG!0�������a��,Y�q�G���Ø!����g�����_Z��n#M�J��H����K&����z�'M�B��I+����1�����j��2q�妙#<���xݫ��ZW�W�;�&3�v�IE���I`cc�\�uU:L�5�~�86�{�j����`��;�3������a�&~���[��IY��Ϲ��?�T��}���]_f�j����IU<僜Z�*��B��'f���نG�V޻몵6.-o��' *)��j�f�8�Q�������e��aj'^���U��A)� Ą���"X*��{�+��Y�L��@��ܲo�b����	��a�A�^B��/v�:�\tϺ�/�] @u�L�z���6 �]��wZI�55�����a��:\y<�ZL�ۮ4��T�嘐|��Q#��͢�RO���c��gxnܨ����ژKGT��̶��vu,��G�>M<���G>�kó�D^�oH˱v�I%վ��-�o���V�k�q���HA3ǫi�؊��%��O����f3�U-��^g~�l�+3���0�П�+j��\&Eo�9W]v�XƎ���K	�H������H�^�=Ɛ�ۚ���g��Xa���U̯Oy1/��}�D5}����#����B�u]�u��m%�Zx�u��Ο�F鼗�>u��:�s��tx����p�����[�J�!��!�c=<Q�z`���a�.^\W��C����y�a��g'ޯf0PA��D�����v���rd�"�㌮J�k�gY݁(¼�f�X�}<F�ߘ�����L0q�Fw�ثZph+R���a���t�@�(��{܉r�X$̛����޾�F'��_�7�N�ԫ�����0�b�	�Q�����m�cK�Ep�����m|F N����z�������Z[�^�� �ICl��	�^�OC�8�M@��93����ZYWJ�\�M�9�O$�ʗ�OC���\�7�?7��`0�&� 
��,u�l���TE�,M��9��j����f��P�����# 9=6U��5�(=�{���G?0fD n�"?��e��|���p�_�����E�'L�eGY-�v���*z�yE�����.,1Y^ԣ�Ƃ&2<�o	���!^͖dh{�Y4+�L����ђ>��`j��_{����#�~]G�E�ryҜ���,�!|E^'�J�A�}�b%Wl���]�Yϊ��{�ġ|��lQ�\��.Mu5MA� ��?qe���K��mm�ޕ�lwĳ)]~x�W�򔸐D���F���1.dgDF�3�����u�s��
��4�(��~nH�<��{ү7����H�!��'F\w� m��yo0g���|zl�[hT�fO��y�7#s_Sy�D�i�Ϛ��Y�dC�Y��d"J<�+Z	4>��ȇU7A%T(u�8U`�xF�gJ��t��T9r��q.�)�#�@߮{ygҴO1�.u����J�s�b�,���*�^��m�x�L���^�_Q`���ғ>������n��*�P�_d� MB���5��尃$��-�m�\��^��˚1��G$RY"*����m��cR�r5����>�F�����������ms��(��|���YS9��{��BRQ#ToX��w���3ȶu[����T����hrF��C�����yf`���Ԝ�y�ӭ�&?0x/�$ ��,���&�������CI�Գ���FN"s�<==�|�#����~&�抋����v_R},�!U�bob&���䑼\�h@�F��v�xw�������$9�U5�v��-C+�Ku�h_Pu�ؾ��k��^يqBF�Q��tK�P�/��һ��'���|Ax49�ƛ�P;6�/c0M^i\�4��i5/ݢ携V���>����6S~+�9��/����t�2�\PGĊ7��<����F�oh����O��d��VҖ�x��cb�g��H<�p8ܠ���]{�h8S��w�.ҧ����Y����ޣ��wܲ� Ld��4޵3��)��0�O	�h������5&F.Q�Kx���.�Ў��/4nO�ԑ�[���n���v#�y��U�Gh&�Y��[�eN�1㚿������p���V�u
�lzr>;z��^��N�4%5N�����]v�B�	(��%�;<0�`�P\&Ҩ��"��DDD����%��¡�2;�y-��'峺_��<�#�W��w,�����nH20L��.@��D�Ueq�#�,\���dA��������/�?_�u�R$}|�أ��j0ʈ;�E/����j�T�c$48����E�:�ڣ��	�3�\�&���\�
[%9�Ӕ�[r����}��	ͫ8$�����t>��V�")������3�.'D���'ۆ��R����{�e #�w5F�ȏ��,߸E��=_���IQ�X�)i*����3m�I��u�Ѩ��7"!�kbu�X�5��}I*t�Ru�gy��غn��99�&���P����"Z�X�I�,ϻ�,q;bN-�/��zn����e�q?^+��[�o���^�lmA�&Q�7�w�\w�n���Y�X�C�@�� @@�?���ͮi���݊�S\JCqi���S ���V�ŵhq�ܵ8	V��]��y�极�C����ڹK~��3'�.�ee���U�B|����*���������1o7KAU�+��Q�SJ��0�g�.�?X����[	�x	^^���q�^�=�z"�
)s�q^�� j~KU��d��Y(�9/��:ܭTX��0�R�E����{�Uj|�Z�LTr�m����Nʹ�ҧ[6n�Tg6�'I�s��_BL���>`�O�o���")n�J��MMH;,}�`�̋Wk1E��EMN�,�e�J�YV���7;AB�x�V��~��==�_Nru��@#�p 1��O�f:��'}�l��TP�
�[��������$Y�I�ϒ�x�ە��A��D�"���ӗ�$UaE�����}v��O�}g«7���H��_�T��GƶZ��^ �ˤN6~��������@��ab�'q~5��D}�.�A�ĳ⮡�XB�w��@����X>�ήK����!���T������g9p:j�;K���Ӑ����g��������wpd�!�ǌ�	8}\�����_m~��(�H���[	&�;*�~ES���ߜ�ߐ�+�t��,Ѵ1o��ꑀ�d[��z��qWsۦ�6�ZYjeȋĪ�zaT�Nw"��W^{Q�Uۛx�dk�U{�<Fh�����PM��N�`��hU�d�_\Gk��(`�gy��A�R��0v6�կ����Ը�h�{tt)AX�%��ws�4�RB��QHK��JR��Y��o"�!F&5drR�v���i��+5�l��C;��/�=MA�D���q�׬"��U���=+r�P��r���2���O��p�j�W(a��3iz��	ڛ'�i^x�8n������D%J�.���)�rR��Xկ����|^���4�O��
��R��M�Дy��K}�N/A롨�ٙ�y��ll�~u��=���J)nx��A�e��?+�XA�#���v�ŮX1��y�z�������ګ����T��cQ��(u���d#	\�ՆT}�j����l�3�b���P���6��ͫOj`�F'�CP���>=��dX.��o��f,̩��&�䴵���o�W�3�_�%���B��	�s�|K/ ���g�M�y�����	�O;i�g�o��j2�c�]5@�<X׮:�66"_^!��h
j��oA�]�z=b<�92 ��nұ��z*���@,�3�#��E#�(N3�]�')�',��w�_%0�Z�>-�뭇��?T����Al�����y�Wf��4PE��G��,yt��,��H����{�ɅL����6b����udKXH�tߧ�X�=/��LOU�w �Mz���[����7��""ˁ{7��A˿b�}�^��C+��>��~���pd��8�ɫ�#����r��Gx����ڰ���a�ƴ�%.����k�%�-՚]w&<�����Iu5i�r��K���j����-�\�n{B���fӢI�F_$�<�NF��aSv7��d���N3cBK �;O�13�_mv��du���i���Pu���R��Gn�ƪ6�ƮnR#��52t5���f\b�q��9/1�o������#_��Px��s�1��������2�sv�9�2�<9MN)�z�{�M#��A�c#��]����ě�?8�V{��F�V���*_�nB������q(��]���g�6�8I�s[�Х���� �`�V��A��N۸\v2\��qZi%(/g ��Yԯz��#g����r����F����lD���[�Й�Jr-c����FC�(�OD��ԅ �2���Q����#7c>]��mo�.>C���l_vP���Se�ǭ#�O�݅�^?`���z����NQw�\�� ��:���O��Q1UG��@�te�U!Ѕ�B'oG�=O��=�9�����7;S�D;�];����������a�Pd�!K�9���m�N/"�[��ZH�'�-�S�^[�x��9������5�����b����������.+Q�7_�6^jv�
���=�-�We��ۄ�e��BM��O�2����_�`��a�*"�;^�y	�Η�f�&ݖؘ}���}V~/���g^�V���e��+�a���:�����L9�(��g.�|��#�g^,b�E�
B�'3/+ս��p�����g�����DG�5"�F��K��!�	[dՓDS�ry��x`4�J�ޫ�ax� �'mS��p�~V�>>��h"V��{_�d�POe��� ��F�HZ�{}������+����� ���s@݀j�g���U1J%��;���{;�����e�J������c�|�	f���"���9o���%�X.WqԃI}�ڇd��o�i�����b�������L���u�$T���~��q6N���JF#��7#�o�}�ȪAG�uԐPݾ��Řd]���O��#��F��<�A�h�?!�jN^��ۋ��g*o��l��熃ߩ`>Gk݌�u^F����ۃ:�����G߶����8�A���q��{�d�H܁���4����, n��U�*5V�"J�M~k�Z38\���AB���H�3�)k��3R���pe���c�2c��~y^��YVň8&�Lˍ5����H���Y	��=��ŵ�؃�V�H[\���k�����f����u��������||!��{*�{{'X�2e��

8/�i���'�D�3 r3�p�tԟ�KԲR�
Ӵ�Q��$C�&!m���Џ�<�^1����~�~�xL�pQ{�M��
�<G��w����[�ʇ��C	!y�H�Y7��wC���S=?�
)m�1�����u*�~F���b�L��A��nF���d,�M:ƭ����ȞL>jk��}�x�,,,�N|�=xS��y��j{�i��+��虑4}�7�Y�as�����+��?_�i����z�̼g"����*�/jhK�XC��;�)��N�B �^��N�A�ښ	"�vu�F�!X�G\,nՏ��������S<{���>��D��1 �c�U!��-DG���[9МJ+(�sk����s�LKG<r
�p<�����Zg)6�j�-Nt~~���
�6�D�J��h�����`*��d�Yxt�}��II��j��6HS���OĉВX'�z 5"@���IBJ*�M4N�+�=�����r�	lzex��:���r4���ٔ.׮�?W�<i	�k�m\�/�q�4`
`ꬷ����x�ڍ 	�̰�N�󋋍L�jwjK�8�7�Z���䊥�%�_d��U	�B)m���~Y.6�(�{�.�f���3?����?�$l�hjl�R@���B�V�R*�����Ŀ�y��iV���)�/L����ȳ���i${C�䄳��7�P�YgV�l�=��;K(x�>l��mӦ%̽�]��}O��$a"לF[WD��M]��)�ݵ�8�����iG���n7��k�gY�9myy�4I��O�L{�o����9:�"r�v�f�~M&薕^�����
�@A����&����71�2 3�I5��sZ�{ā�9kS��O���xm�K���j�T�u���9�0�F���Dp̄��<mH���C�9`mwiCؕ�6��{fc��k�%�B�\Xc�O��% 
]����魆l��)
�T/K�Zv7���1E�>E���6��9Η��y����ڔ��T����u�ZM��P:�������z�8�^tJ�Ȏz�(2Xj�����Q�0�BP�� �d���ܸ舋�C�����[���efy�1��0�/�8��aO\��V���ʐL�&ǜ'�.)5��n��h�bS�);�ro\������ۘm�� �A��E}pҕ�R�ep�v7~+s+n��E�����Ĕᖮg\�[�>ΩgKp�(�nk��4?L	�aw���RɎ����~�A����[v��o������)��qωe#K>��T#��
u��u$˫��޳IG�&T��_u�����y�A�~ü�k֐�ĸ���Ĕ�s�tZHk����2�����f;���Aۭ�b��\��eX<	l�X��6�e�����S�Hl��W����Z�G��m}6 �X�5���x�h��m�DT��� �>��9����.*N�;V'���b#�p%+kT� %��I�Ml�[gD�&ݜA._���:��O�{~�˥L��<��f���t�~�e�%�6�Jq����zҘ�lW����m��U�Ɨ����jS���S���ҋdۺ�\��)Sᨂ�6L�|
��'�N���}�r�sX���,���E;p�|��F��P�B���[���B �^��M�I`�ː�e%W�i���ճ5�Gx8�A�0�	z�S��L륚�	G���e�zxԓi�~�CV���E#6���ۗ�N&�6�Z.s��s���p�|u�_p"�$nUV��r�w*��Wow��m�%�Y����˴!�k*;	��O�Lټ��5i[�dj���*<��fKQ¾:�ZC\��� %����C�i�| ���"������Y
���t���(2��?.��k 	`���ƿ^��Z+�����R�fk�?��no��ı���]G�F0�D�A�ƴ�~�}|����|���٩�ZY���cԊ�JU1�'�[��13d�U�vY��^��>@K�\L�m�c��h��K�<��I/�3~��4B��'�Z�<��1�;�7;����n��cuC����L�cy;w��]�γuM�~�Dv��Dni�#���W+�o��.�m���oO-˗Q۷"czs���گ�311r���Ai_�c����I�j^c�D����`aqg�0Q)茍�`�ض�(�l�}��Ôp`<�aHP;]Rg�]��lx�����#�k�J�5�4�"2NHU�?�Ѫ�U_��b^Ub�*���S?�N?��v�r��G!�͍LL������D۾����^%t�"�� �'R5R�S�Bf�;��^�s�}>Y�����41����6"����-�dU:�ǝ���@<�'���6M�OY�_k�e�(��
��ǰ�T���@���C> JD9�}�����N���z��gJ�%W�r�~�&A��:�xd���!�i��'���V'F�f��S�/x�O+u���*/�?7��|�T�-�d#���H'��v�ګ��R{�Tm�l�@ʫ<(��8<��9���=�ݞ��8q(�T����M9e�����!W�7��8i�#fǃ�6�{~a�Y��"6�K�ΕW}2y��9B�al�Pp�nΧW�R�4����[�����f��Nl�}�~�eOm-_���6�t�(�R�~��}I!��;vNU���߂\���őD�{�@���uM��i��-e�߳�����1Ѝ���ظ�;S���GJ����Q��K�r����9�ҝ�e.$ѓ�U)qp��4�vN%<��,)�"������h�L%��uz7y�m��`�`�_C�f^b���Fm'�PG�gD�B���9�)��ׂB߻F����P`\N�ާŵ�d��}&�D�/c��פ�dk.O=�8��Q/�|V�WJ=%a���UJ��o���������\�k���B �Ͽ�Z=��"��i��0	Uuu�$E3䆜}���,�S�E��n�\9*Ȯ�ҩ&�$�ʎ0Ɯ�SW�,D�lv/<�����Z0譊���z��LH�q0S͌�?���������f����z����bv����L)1��h˫l�	�V�����\).��3��r�q�W�6ږ)h�?�ʿ���i�l^��T�v���w�m=}�}�i��Bhi��X`l�M(w�Ӎ*y1�4��Ŷ"@���#>Iɸ�#�:�������6_S��c)z��f��/���<��ue���&.bEYY kX�_+3ee�v���P��s��� �{�I�m.)^���f"ޜ�א@e���� r�6���b�ۣ��W�"�c*�k�|D���U�۵�TB��t��+���i����,^��f(�ߥV��6�\>��
��d�?�	[XV.�O`�[GDF�\�� �����71�����{o�٧Fجb����̷�/#�8aevi>r��vN�=��k�B����7DCz�?���pc>�����W��
K?L�����t����O�ǲ�'���/���\�-�0�)���-:X�;ݹT�t�~��,�f�q$�m��B�D���/�R/�������[����%���V��L�i0l�#�@�㰕@��� h�_�������va����YEs��ʁA+�K'�>+[BT��rΏ�/2�eH����2x0xڵ���I���S+�Ab�eDp���1�]š7&�'Ϥ��}��(�Iʱ������fܮ- �Iw�)����'ө=�){=�nD����x���ɼ|ʷᚍv-j����Ck�hu��@�i����F��ْK�O��a�[��['��Z��r�������#~)޹OߛtW��J�+h0�1��Fޠ}�¥��z���K���sK$�*�Xtc5{�o��qew���g�}�HJ�
����(�.ϯ^��,�L��x�5t����,<<��J|gmPN�
8��w����.�@#s*�%b����B?�~�30��Ya[����Ѡ$3�l�E�/;��O�J��F&�Y6F��k9�-НR_X�+6@�b���;y�Yμu)[ŌVP~(��ݣ@I��<�HA�I��'*>n��iH��-Iv�g�!����1=�S����O҃vS]����hy[����DR�R��ˑ�6��c5�ӯ�1�|�H�yFi��F�^�p'	�'��Q�j�.;4��bn9����n2����� E���׍�Q�2��g">:�#H�KKli����/+�hE���B��s\����1	7���Me	���1vx�^��?���X�0}�2�TJO����B�[�f�Q�6_��ч�Ē���Vnn�2Sw`���n�b	'wl\��U6j����6�C���K�tC1b��"�?���f\2���r�9��dL��%�+�l�FQr'��q�OQ�~й��s�z~g�m�v����)Ns���?����<R �m�qCbʧ9�}��#R@W�٬��VQ��*6�[a�<\,��M�V�R���vX�\{V���ɍ��@X"aƟ�A备 �Iaq�t'5��b[���@��P�-���ܠ����7q����	�o9�}^�O+\0=
H���s��qs��|�s�ы�6p]�I����'����V��G�VR[�v�OI�����|52X�b��o���]�U��̄)}�1�'�6���5�W���2�vÛ�a�07�T���ƶD�^��ߋT��yF�5�(�T��m�����͈�v�)���HխA�o�U|`3J�`O4G�˻�~���.%"���]��7��^������X=��;в���oq�f�3��2��}p���(~��	��*�Rּ숈Ӣ.
?P��ԫ�Xf�*�U·�W��Ry$���昕�L�_ ��Bg���t�f���bײ|}�����E�(��aqܳ��+��@�?7�e�dRe�j�zٴ#vJ͎��)30�$X��!?�'��u=cod_C�D8��f8�����O��wlmm�q���lj�e'��K ��v���=�2��b��Y�=�a�p�BG?��0�|�lw��R�g��`CD��}�|v]���-���O�(�"�k>�Cr�
�=gzM���P�NT���<�3�l*ƀ!�R��,�c��t)G�)W�����ץ|�f�C����4���pό(q����8��\�wZ���4��sF����p���gf�R7�M���>�s�AE�a-�q�������D���Ueړ���~zJad ����W"�`�,��+ ����T��l��i7VJ��?��:��Yn�( �S�0�k�K�os�}�\;7&'�=�:��:��6�����
F��3�
��QG�{</=9���'�c!.!֕Os���h��M��p�E������ԥ����!���jS?�LG�@���;���,�a9\��M�Ç�'Zp;�g[�z��I��q8���E�� �qXb�K�/��<$�\<���֖$��¸J����+�:�G�k�N)qS
�秃(���8�͐˭gX�\��GC&`C���8��S�Q��F�1�A���8�;,VW�4�]=4絺^.&�8��X�樏��Wk��{e����΄����=xA|���������QtT�A����ʊ�����Jh�X���kv��{����'�i��c�H�'���9 ��,��3��¶<LNJ��Z����}�O�B��j������F�1��͠n"{V�V��y�?N�j��1ï��UT��>�ꘗ���i���k�л��āI��6��+D]Rn����%X1���%*���qcIa��6i��� #u[�F���$d�g�(.f�$�����@
K��'�O#�	����v2�GO꽯��7UoC�������ߌ���X~7��憨5�Y�2)�&�4P
�VM$~�b�`HB�:%j(c$��k����xbqU�&�q���N�}ԝ|��.�;�e6u�~���`��?[K�x?>:H�*�Z5�M~z�3
�q�u}�f�wn���2�sh�D��D���?c1{�}����D�=H0�]�%���]Z���ᴃ�c��"�	B�=�b�?�'�ž>ݚ>q��IK~�������M�1�B!�������[�]��m��lf<؞<H�N{ZX��x
B��t1�dD2�\�7��7��$2�� ê���E��!dlr�����)G#c�(4-���8=wh��$�B��6�}�b�{�S��oh��x\8��
htd��n�su�W0�b�U<���/�? uk��r�vR"
\�7�u����˝+>6Tk�P�� z)����ӯR��"i�(��V�S�"���f�k1���p%���������]��l���Y9�j/�U�_m��Sa�eqH��ث���d' ?�)/��a�����f�(�N��Ћe�!D�哊4���u� NrYefX�%N����I8�*��k����/�6D�Md�̟��.�n��Mp��8�>���4`����p�r?gY4���Z�V����^��p;���tDb�ͤw�׮ۊ. h�EW��I���7��Bs�:�d��}'�W�Ќ��2k)�����`��Ǻ��x@L��/L����X�"@as.��õNj�6�;͖����t��s��?����眰&��&p��̄:}���,3��Ӡ�<��[��
�T�{�u�ZQ]}�V���J��� T�:� ��]�:�q��%܆Fr��_�����:ϋ�)��4��_�{���(��Š�y}̟@���v�V	��LA��!�H����P�M)0��H*�d�9֩��S'���Ki] � dCV��"AjK�G���ʚ�GZ�s�e8��H~ZDO�P3^�݅�
>�Bs�Q��O�'���ѳ��;w�ąLЪ+�\�P�?��
�����a�)��������ɷH�Q6�ZL���n��T���d/��}���u0��k!Vw{nx�'�$�(ܳf��y\`�(���#sÅ��::C���/}ahHw�9u����!p�ehs��=�_������$��7H�|
�s��ya�W �&}�M!���]�L�qȿE�b:a:i�G�x5X�w����H����Γ���r���p���ǈ�V���0D:�ͻ�jvw	��X�W[�Z4�O�擾����N���U�e�w�cW1�pk�3���4�M4Ņ4�:&��ƛXAl�lHL{IX�[��1 ��Z��µ&}��a�<���^�C��p�#Ϩ��}�Iu�˕J<���)��'���Q�(�+6�4��#<Bx�`�|Dpld�&�i����I�]7}�V��}�@��xA�_ӳ�>�+�m�l�2T#ny�6������f�;௛�"~I�%���� �[���S��aqhh��K�!41�^-���d�ŉ+��>�5�����q�a�0�R ���f�z���ƹ�NW�<���p��	�{i��<�6��s0�3����CG~w��^���N�k�0��K�>��z��#�ں=�A|����d	��@+�����vd経��j$۶��ESd���ZI�g��7��:学>J�_a�zp)�'ڱ�T�T{-J8��X._���UD�]���ʿu�i��Z��Ia~O��E�?�\F�Lr����޶�d�67�^f�y�Z�ܶ2�����}:/�\7�[':::4�� g���p�9ﰁ��o���Jp9'Q��?���Ԧh�'#�ku��j?\�s��^α4�Y�Fv��9�4'�� =/s�9�w�z�Em���}  P�
3�'4�\���r�	19,��/0X�ʁ,g{ReNrV��%6)~ءG$�8G+������rY��$."HJ��E�+����py��ߊzQK�A�6#��@7���,�F�,���R���վǇ����[փ�je,�=���z���87�(�I�T�������A��̍�0�,�J��_5�	��Y�ݧ~"9匘���0�Z[fs������a�$+��[LІF��/(��i�E�ǝ�kymZ�i�Fl���7k~��@�w�+���9��x�utt�õ��w��+E�u���x���<��X���#�|}q"���E ����g��%זTYj�I�wS�?�2X����U�*˺o�6`����[�lIX(�fOl�ÄE�� �,���7h9E96e޳pǜW�M�ө�KOD-b�%y2�MF�
��)��
�����Or�R���J�vu��A��f��)�/�3Լ[Ϯ�W��@W����S�5�ȱ��$F�i��C��&´hG��%�6ȂP�S�z6���D��`��*�-��-�o�c_Ӯ�M˛X����g�cW�R�Y!��`��{\U�2ȁ�c�!=/{`e��_�MŇ����P%�WN�P=��Y!�˅:�Q��
*9���k������#�8ǜ�$B$̝ &g�s6�%jq�i���WBب%u����A�Q�I�Ǜt��f*A��o�E��xy�bM�:o�kx5�;>�* �/�_�|i�ܹ��ZC�X���<þ��[I�C˵��@���.�F�5Q�#ݼ���>`@���EA�g���y�}�solXm����FJ���js"�Ε�P;�E͑\Ϧu�L�]��u�A��L�-�̇7癡_{[���������H1�V�]�k����Rs�g���8���m��GR��A�x���-3��\?��XK4ti{���]o���'�IkI�c&��?f��IL�����^+�8ތ��c~5&�4�Gl�%�ǃX��[9Xzh6�gd���%��j�/(���1��+�A4�թ`E�@�	-W֜S`��� s䄿~�B����+T�]��y��"�c�aR?dQ� ,��)�:Ơ!�Ѵ�� ��,�)6�}�{H��2nje��~o=�W_�Nj��׈ti�e��A3��%s�<��G
!T�{ŏ����hd��Y=0A�P�� 3������%^Odl!J/Ϝ6	���L��Ac%��
�&$Σ� �|4D&���հYZZ�/���@� :3�D���]���޿���I�������=%����G%���Kz?/���E��$�eKE]>*o���OH�A �8�t�IX��e�ʖYe������A��F^ꇻ�_���6��@����E�=v�λU��Yޓ�	�[3�Q�q��$�Q���3����lBA����J��ׄlON/cq�\��@�2�0p�S����y�> y!�Hu��q�������������U�,˅����T?�Z�	�� ��Z�ɡAߓ4
�{N�7��=�q��i<��r=�G�Xi,_u)ι�x�/�6�]~A�ē��!4��F�A1�Ft�r� KFc��Ɣ�Hܵ!+�b���/)��3{��K��6�L�s%��R"%]�GJ�y_��������_�(�sW�q��u�c�� ��3�v��B�E�m�n���`-��
�;+`����d"��fQ���9YcL�ĽF���^-G��U����B_�����h�;�Y����0�*�����b{S_��S�z�3j/���A�,4��ϕ��REƆ�ꤤ��j���w/�����ǩ�Q��
͈��*;T��J�Q�b��]˔����+@��f�par���Pr�Z���f?I�Nϔ��$p`�ދ���F>��⤍���q���2���ϟ/�np�DfŰ�3�M�I��B���/��v���v�Q���R޲�i�`�}�S�	�K	zC����[+#`��y�j�$A�*�ưn+G44�:�@~zzz>�f�Hi~�{Ǚ%�!Tz/v�i�I!�o%���<���ķ�����5F�n~uh*�6S)�]��_Uʂ\ԅA��ĕ�.��V���@*��G���I�w���/Lb����9��9��������y/�:ti�sV	��mQK.4!��A�),�ִx�[�msy�Q�7B��?rz���>>7G���ؑ���xn��B�Ecw.�d�${�*�ڍiW�^V�KU��Ta��r�E&)��p9ʲa��K	���x��-�L��@Xls0,���V�����"�湤�ԁL+�)w���q���t"(���2�ȋ�ܥ�Zy�ݦ.�*PS�Y�{E0�G�@���y�)��4�`����iB�ɜhS����)�������/�捉ؠ�/	7=�huPpJ�+rM�z�[ЛC�j��'��l+"IT���w�'�-�W�-���eT�����[AQ�#+~�u���7w��+oX;��*�2L±�Ɵwu �ް`a�n��`�Q1��j�v���w�����tS���%�����aq��aS[�wv�N��4|����r��%W�7��X�R��,���-��@w��;|��b��ҡ���b�B�E���b�K&��y7AFs�~������77&_��zu�mrqb����;�wi�r�e1N�3a���I���\�5@"�!��QW�"	�=]X7r�9�|�����,|��A� ��p��33������<'�M�t�W�*�t�:X d��E�q������+�n���� 2����^Y0~Ju����?��/l���Y�ƥ�l�G��d��.uTV��*K�.;�}��p�&���[vk��&��ps%����z�?��ٹ%h�ݣywN:<�N��h������ia�/��A��ỳ�Z:UTT�p�"���f�n4�F���e��!_�KC	T�c�N���"��>��1�R.� ���T+^�:y�/H|lKtP��?H9��d{��:2%^�3z��z�%o�#���ZG��W�&����d����/�Sj��bZr�p�S�ؾ�0:)��� ��{ҙt�6x��<�=�]c*ĥTB �n�������t��]�8y �����qe�A��7�LP�	���P��zql$\� @���חY8)|����Ȁ|Q�C{��G��e���� Gr�y;PP���߮]�l"���Z�b��}~'��d/�%k���܂�wj��m,�钸���sޙ�D�2t�;�K8��/���Y���Tze �b0���+� �Ϡ�=����C���KEv�����x�a��Kŉ��0��ǱF��?���F�<3���2R�_Ah�BA;y����+���?ի��F-�2�!�Ï��f��Uܤ��/>� U�{QT�ܡ�qdٝK/9�U�3�
V�N��ɥ�7�y�c=��0"�?����C#9����ӄ��n�	��>?����2��N9Ed��?�X��(���ѐ79��F��IFӋ�ȦN��JU��Þ3��E9O����"�;-)q�}R�x�ʭ���m?�t&�̷êO0��כ>ɿ�<������تb������� ~)wD�2�1&W������9~�{_2�Z�@z.W+��3v̌�U,��[�c�tX�j/��w���.K����ҳ'��b��p	���Hd�F���9���@�z�Y9c	�����V\�$<۠k+�k6�sAFv\����������C��t����q܋-
<$Of� �1�ڴ*�u��V�������߈�r�{%��O��%�7/%	`T��9|����+��G�
ı��SsQoph�T��5>x�Eo��Yԡ� 2Mpf�X^��� e^�А�K-�È��D4�B��_l=Gz�t�����~���ʿ���U<�t	��tԎ�F*���C<�ŵAd�N��S&!1CW��x�G�wF���0������cP?6.��Ǖ�[����p�7��ޚ��&���Nm�)x���
�j\vΖ��ݙ��C.D 7B$�8C�^+�Vi�>EbH�f�[oYZ�V�#�L���s����W�����إfg�xo/ZIi)�T�cݛ�o��cB<YtCZr֣��'7�k@Q�g��Ѫ1� ��Ԃ�h��8L�U?�@�8?Ĭ�)��㆏R��5etB��<��M�^��cfj5�z�N�ww���ju�qR�0LS�P|���A�!�x��n�2��=�(p]�_?���=����4�)�t�l�$�u������{o9i�cU�:uV���Ŧ���.\7� v��ٸ�XP�)���lH��ޜ�����y��Z{_G�X�5�:(�Ғ��S����}@�̶�ٚл�1*p�ճ64A�0���B�"S:�s{+�t؛SkDk�@:�j���4���l)�4c���a8dXޟ��<���سŽ�~��G�vw��M<�I��eiw`w��(31(9s
����s����(������XѾቃ��l{��Rn�\/RG�Yc�[ϐ����n���\澴4�ޓ���LRx˱���F��,�u���U>:���|!H���?�.躽T���EѰ���"f�L�n�C�,-FU��O��n����^r*�pL��7�@T�<2�>3՞u�	�ج�wZwgm�&��]7�v��3�y%����7��X1��rNm*��լ����M�KMD�t�0��}�+���$.�z��P.Wu%� qzɲ>��m�R�c��Н����~��മb�a�i�݌c�.�y6;���-*!�A֦C�g_��p��@����4��8�z3���V+�[n�������h��Rm��`!�Z
���.$�W�[T��Mr��/w�*G �gF�4ۈ��8jJۓ���\nPݥ�rMQ��+>5��wڵ��v��R�>m[�Vf���h��w�'_�����{�y^�<���������$�k�~_��;�mt��>��H��H��e��?��SP����Xw�R8�PЫ�~�Lg��}B�C7#8�M���U�b���V�¬i��D�B�{i�4:uP���Uׂ���R��<�J"���/���E��a6��f��#A��(鱐%MH��Ĭ�E��ó?ۮ�*9�P��կ\:ux+s�C�X���T�W`;��sN��'�R q��hv�1��8�~Dd��q?*���Ӎ5��j�+�4Ҵ�"/-2�F�X�5�)c�X�S0�
/�i�g�=s�*A��V���zNj~��.а�E�[�~���ܦ��޲@^��\=����u�cqS�����x����,c��q�;C|�!�-f�N8QbDy+���h|�I�}e��=#�)?�"Y��v�@�ʓ��'/�E�|�Ghʏ�+v�dM����$���Z�C�m���X߂H�";]��j�����ȝ��.��&�;��O9�W�Lۅ(�vK���l|�0܎#���g]dE(ɕq�&�̶��-�6[��`��3��;��2�g��&U�&qSBg���r��;��m�9��;��8O�aP�C?;�`���+�-�zӬ+[��!qI�8)��s3k+��7T�WWV�)��+������4�[��7�]��6�o�J:-�N���@��,�M��UѱnI��]��P���g�cx���=�K�=��E���E� �m��%����"��8�9��kf�+������֓�;���?�L 
8�ŕ�҅��V�H�����H�����e�܉L3���T R��Gl9;*�@�����ĩ2����"��A8`�eH��0�oE��|� �|�H�E��S�MjK�7��d��P>/ ^��:WN�K���������Iim=�&��Z�(�qt�In�ڕ"F�m6�Ra/9�����͚d�]{{���`��v�}PIB+���[#��4[��A�EZ�U�A��!����>^v�W����lې���!����s���G�ru��N=��>T;�m=����K
U?�J�0��-�HLyG'�,�.�F�5{�]b�o]!�(��%�v(�e7�W�W�����5>�͔WN[�����R�&��:_{����TǍ~�7LUL�, ���������֡���|"H��j5��R��m�:e{-�c���P�%9w�y"�:)M��ra��U&�PO`��\��^4�[g�O���ȼ�����C�ɹ�Y}B�'��ƦI��ձX���õ��q�7����l�����	�? �j8?Ĕ<�{X�q�\:Y8HR������� Y&�i�N�̅��p�8��/@�&)p���V\C&�Cdl�wM� �V���I`:7A�-*��1�����aM~�� �"H"%-- �0P�S@iҍ��(	�����56�cҌn�F����|��ϵ����y����_��<�9g��n۠ϛy���G�M����j�ӇY���R>�����u�z� 7.� �[�z�9�� �L}â^<�}�޷*�g�l=�Cdu_�F�E	��4�]{# ]L��/�
2�D�-�e5��l���x�g�JzN���V.%�T���5�G|9�� �%�#� �fI��yxe��{�����~�����Mءl���������_��|�N�;��^s�WI��(�[��ģ���շ��*� \;�|�v�?9��1J�f�s�?K�8`�ĢMZJ�򬨣���B���f:��w��ּ��o��~��{�ڟ�g�A�ݼKݛ�?:��z�۶VS7�`��sj��8U�邒.^�H��(xq�V�@yyz�m�-�I)�A,ǈ��
vA�>������[;Rj��/��鍫�x���7��'I�Y���1��˂e4�yPږ�v���a�����{���i9-\�J��n'�{�����.��˷��	4�ˠ�HJ�=Xc�%��ɭ��m��ݍ6S�Ԛ(�~�O��������u�(��x��S��}���3LDݳ��p!�*�;+��	�N�u/+t��'��&~-�Kɽ�GZC�p��E��	���	h�)��1c�:�u�:I(#sz�<�M���x���Fz$��2f�>���G���X.��� h�/d�#ZT�l+�;�22y�I�'�Cd�m�g����{E�|��=nq����z��ѫ��mC�HD���;L:/�` _�n�*�9XÂM!ȅq��0�ĐK�t�=8�\)�ޓ���?���J�}�@��˱ǖ����5��h�,:���럒}s����u$�u��}]��摵�`Q#�ȓg*��ۛ�*%�������Z�!G9����� ��D�I�@��NLB������C������z����-�0iǈ�4�g//��Z�?LEz���
9��#��'��a��7��L�5ng�_{uC���ւ�[C��W�i/.O��=���(��J�h��Oz�H;�3,��NE|�Mi�d\�;��~�:/�5��	�E=�.-P[`9qN�W �8=n>prT�ϸ�:�����9��W��o	y��Y�t�qT��߂�V���0R��Xn!���ָR�B���r�.Jw��^�gcI l�N�4#>}=e��r��k���:4���W�0>�^p͡D�3�Ӑ�'!:\�XbkŻzjh��G7����,�E9��ID~�,�=/{�A6U�����7{cz����0 ���¡�,@R)q���\U>Jl|�����I~s�-s'8*�;n�n_�s�}U��ѳnc�w�r�ҵ.�<�$Ty�x[�o�} Sg&b7L\��dXp��.���
�i���]U�?e3���oC
��% a�<+5�j/r�O�=�2���ѥ�yr�}��%����&
����MY:T9��n��T��d��og��Q�5�6�W̌ח5���M�*�OB���]V}m�LE�B�����Q�L^���j⋼9l��Y�Pwe?U���I��f�4|��5����WeJ���l2e��I3�g�z0��r��^K.E�������q
Ċ^DR}�M��܂�Yk�%�_��uKىrQ)����[Q�B�q���Ie����/x�{$�t��z�az^R��E[!9�������y�a	݇�{��E����a�Z\���Ř����k߿��?�v�ͻmd�=�}���n$'��S�T��դz���Z������
���E{&�>%j�g����������o-@�R��j\�HJ	�:�I�qљ�S���QҖ�!/��ǥ�T��S��Ý+�L���1�}�����3��n���kF��[�g��������D/��-DD��)�{F*�e��=�%����7l�8�*�HY(yj�1�$igw�sZq�0_���3 4� ���ο�������8��h��P��6��H	�H�[br��7�����N~G9	�-N+^ H�8�����1D�l��D����X���囈Юo���Ogr*�ˣ�e*i�M��o�sC)ԧb�]��C-�m �%�Y�z�fD�g���3�����K��^���=Vs�"����\��u��1��}9c/�[��N�z��X�?�eF���]�nF��>�UkY4�9�gψ�ˈ�YV�����ڸ݋t�ͷlI���}J���gMM�8���.�|x?��Y�힟���k�憊U�qC���A$��ϰGֳ= �e�+��i��ހJ�2,��ac�ޖ� ��ė������'�=��_{HJ˶߇x�o<���U�|B��y���j,���ݲ�`�T��H(�n8�V�&[qdx�S��\|��s����w�G�-��ϮL�yx�y�d	�%�w���s�)tzo�H��͹?���6���F�[�$$~,�~̴� 
�.��Tj�n�,���`�ѲZ�7��"�CO�:f$�����D�����-���d�����'��⧎���m�i=a*}T���o��'�L�	����w�0c�rRN?)���b�G)�&���3�]�3��,���9yZ$�����KjU�a�w���t22�V��F2����l�9_�{�͠�i�J"d,[(i��YfS_d�N�sui�̬��^κșs�}��SPa5-p ^�I�s�[9�C㭶P�數zvw�����=�l0�{�0�KCbr�l�	�����j��ì��*�(���&��\N��8���� �	��>��L>h��"��RIE�i?�;����6p�gQ2]x�J��N�($�'陙vo�5p��#�
��Q3r�Ch���2�QU��W���vf�:V�����'��/�j;°�e[p�^��P� 7d"���ǲ���sxPis��%�絷���ˍ;ɲTQw���8���^�Ϯ����w�Ҽe�w�-���sw@�?�`̷�ZI��j�i��$���D/4X�FkfW\O̡86�ԬKЄ)
)`�q
�e�B��4�}Ob�e�;|[��G��Յm�aq�g�tPDGb6�05���)U	��.+���!G��5���O�=<B�Y�O�mm�@�Q�ȁ7�����]�z<;	ųLBS�k�$�Ԗ��?x�[�YcF��_Y��o鐜�M��q��څ:Q�J3i��p�~qJ�Y�;���@����K�L�#��S���|�h�����d������F�zA2㊔h�}br &`�������L�����W�x$fL�f��/�ǌ���S���s�%���+ �/�����Xc}k�R��*&���F����z��g����zc?��)��.Dkh��� 8Uj����#^������h���q�-��&���?�,�s�>�o�,xI��e���is��̦""4ݳDz{�H��~te�\rY/#Pݴn�5�>�u[T��+>Y�W�e7'�7REI��H�r�sF�5z�=�ْ��nw�<��<C/�6�Gb��_�e�ܴC�.�[���
4�ɥ�T��]�Y�d����А��0�9PG2	C���̑m���N\̞Ϣ�^���K}��w|�t��U�D�{�M~5��V|$�ɴ���*R�W�Dk�ݚ)�&��<�:n#�����z���B�PS��J��G.��'����x� �=�Pm����x���5.�v�l���l��(�|g1�l���̅�.�.�������L��խ��ݚ2�1,	!��l��!&<³��"_G��k%_�9vN��1��z���.�oc�x)Έ�6ņ����]�}�6,^�8u�~�|���X�e�
cJ}��-_����ߗ�뻗�;�R�[ 2��q��2-���'7[�9	�c3N6e&	�s�i˲��S6�m�!wM�.�aB�Rt�O�R��[T�L�\3��m͇l�����E�n��T�z�2���#�?�3�so��I^��]jFj������¾~�����h9�V˅�n��BHm���F�dn��^!;E1'jkm tR�ߦ�"#�S����zC�@�����ȧ���ֽ���K������m�o�aDYc,�O�؆�G>y�y�L��h�A!�B�0�aFT�eS
F�1GӤ���'U��@/{�<?.��te���8��gJ�Y�s�z���1�l��$�;�QY[��_LN��.� ˖�Z&Gu���:�pR�S��ޅu�犜��'m�ݏ���g�$#���""�b&�/f�$���[�r�f�j<��x) p�d���ϛ�,���S[��"v���9D���χ�,�I�m����R���U��B� P�oF�U�3�}M:[��)2��d�O9Xx掭��� '�t
�����S{� �{L\L)��o�)"`���i?+��z�v���(<6>��ώ��-��B�G�/�^�џV���yTS�Jͷf��T�pU������� ����	o�	�V>x�/�����*#�ڝ5:P'=���]�ݖ�N%߳�#^kA����xT����!��?��-F��r��G���ޖ~��̙�)UX���IV:V����tS��y��\���>L��Z��݋�vgv��H�����9,6FW�U�6�/�v辞�y��ަ��m��/�ʽ�8f��1x)�+f�?쒗i������wy���kJ_��� �3�*��Y���^�z+�]fa�D�\x�?��(�y���������ß���+PϢ��nߞ �̈́�`FJ��ֶ��4*uJR��u��x~踶*�+�~��k�/5��Z�8o���<������k�!�H�N���������E�-��=[c�7t��=�ǝ<���������gW��c�Ԗ���D���Y��G�E�DF���7��Fy"��ワ�%�kL�&�1r"!�f)e��ǋ������co^x�e,��	+�.���sI������s��~��E�-y�\A	mFM�����M��&�vn�}I�w����r൥�]U���{��.�"R�HO���兔���S��r��&��/m�0�e'y���;�<0�<�I��VW���$F�,��!���^��F͙N|�̶�.���o���s��&�ϙ���M PjH���B;�������cpl���U�;�*�����tfͩjn�U��ڗ@F���{D�AW��#$���o�$F*���Pi9r^�.�=�	/��u?���{��qZ�o�s5_޸�}�fh��#�
yߦ}� ��Nt�Zs]���4�,�u_A�:�hR�'�j8����<��.�c�l 

�¶m�ͥ�T7N [0�cE�GU��UV�ќ����d(~APl�l�Oc79�f�rp~27�����m?p�������z,����sة���xʽ5�n�ߴ��	�2�0��砽�(��ʐ-�V�� ����޽`b��;�])�z~drhh(cWW���K[��k�'�p���g��;n[�N�w0� �'UpO�����ĕ��W���d��^f�Iwn���+������ey�����z
��w�n^�bK�r�s�"���W�B��x�'}Rٳ�&��/�(�}��t'���4)���Qg)ה�P�ѷ&��������Y��Qzڨ�ٿ����j�O/xy��Q܈��(�Y0��ݠݚqW�y�j4R��6_��2-���3v �9;{C��|ܯx˙��������{Ny��x��6&��:5�A�;�w��?o�lu�V�Rb����P�����M�Gwg���:�r��u�fy���S5Dh�J��E�m����o 1 %󺙏�h�G/)m�l���#�]f�<4���[�G
�Q�ڑrMe��<FNe���Ĝnx�>��^{�d,wz���W���UĘE{����f�7�߯d2)�4�����Uv�Q��h�1E<�a����W�	�[~Y�=L1�}m:WB�H=�+��%#�ss�S�)w���[����m}�<yl����`��[ie&�0O}Uzq@w�f�SCWdсc1�k��*b3�n�S[
�^��P�Rz�Jfǲ&".�Tȷ�Y�B]��f�f�Q�,�bhRM��o䋙ἤ_��n�o =!�R ����MAb�
$��0r����? 9����<Cwg�+7+�2ԥ�GɵF�׾Yvηb��#�Ut���dk%*?;��k2i���JE��d�=����S�[�\�v�;c��N�%/��V\,<�Ҳ��< �߾�m����2�ڶ�Z���kɐ�^&ܬ8��]~hχMXG�hL���W��ߩ�@xZ������Ϟ�����Px������BKR$�U@�~/�`]��Û�$e9b`����d�25e�&�L
Ƃ�Xh�����3�_(P���u��,_%�d���i'�M�k��RP��:��DS�����툰Pb����ßO�8�iv�䃻��M>_$*��5�_)͍9	NW{W�[iox�G�7KEZ��=ܡCo�
2H�����ޜ 0x/�tϯd��(1:������d+(�A��f�e��
x����L��m�ܳy��D���������0P?wn:<��c�r�Sc�.lr��=]�.b�M���Mϻ3""`%�>"p�&�f�F��nR�<�k����*V��ms���>��\L�ܑ6�n��p�gR��*�G|K�aJ�����;X�}���K��#���M��<gY:h��v�2%Z�T�#vgE��٭��k �t:��;�_䖑g�4�9:�����n��q�C�U�v�;X֬�!:��r��JD�~�l6K����kF��V�^u����T��B��F,Ssh�3�-�YT����/~��ސ��"m�=���w�a�ڣ֬��Yc�Z>�� ��}�r0��L������J^���)C)�s�_�r��Զ��p'1QX%�!��)QR�2�Fޫ�E��Z��$b�1��W�t�E.�"��=�(��[o���@ �%�p�a]E��̫l�m]��I�T��]����O�Sx]d [��x�b�>�JP�"��h��tP?���1Ҧ��lE^��(����o5*�~�&���w�m��m��0)�E\1�}$K��C��#(u����J����gd)��;p~�t
ٹV>|�#�����=g��$0�,��#l�z?�㒝�նb�������(Sz׻�'�����˂r�\/����LH�0�����=9��]�aO�/��tn�J6|O�׳�"`C���KF-��M��|e����5��]��	������1?�]qD��iTu����S���?��@%<���x�m�%~�bB���-��Z*��	��^�s�د�f���m�m7���=Y|���h�׵I�4�7�ѥE�H��aR��f�*$b�������Nv�-��3y�`S�AD���/i#��S�����\��w�3E�pj
����Qæ}y��NN��d���Zz�~��ސ�߼�wې'�j{cV-F�c�O�mX��o6�?iw���k�:P@#��d��1��۴�
�m�x�>$J�-�Z^52S�ߵf�-�P�ճ��D����������cUx�6�k�K�+/�t�d��W�:�^':�{�j6�>���v2�;�x:��
DԪ}.�M�y�@�:�QQ�����Vtmv�w�e���л��}�=�5��R�����9dS�������IEj�d?p��w�=�cQ#���gW�k�4�;���[��ƽ�%E�or�[�k�K[�.&����{��ҵ�H{���������ly2�k�(dv���	JKC�����]j�k,ң��պ���X�,�hH���������̓�mz'�t㹮=�`k�����|:N�|r>�C����7 %3�z����{�QT��T��w�O[W� �ڰ������R=����(9���§�M�DK(a��h�qZ�A�����	@hL����vd���Vћ�ƛ&b�0����>��'zbh�K(���s���Et�m"�ɨ��կ�QJ���XsZ�_w��-j�O��'k�e'�ss��ÜQhC��O�'���}D�A�@-|���K���ڸ^�>����	�o<W�n;�7i�|�5�'_3J�>��.`�9����yL��uL�B�{�RlB�s$�@b+����NNZ�� 2db�qJ쀯���ƃ���	� x�+q�>`4�{��ǡ�%m���C��/;8�_�G�]aE^�t��ж����]ܮ��w���������+���#8��P֣�/O�����{��\D6@u�bꕖPmd��q�%�����S�}��)*@�0#G�4:� OQ�:9��ν�b�Z/
i��<f�����!����m�+��Q����}~�)�ci���ޠ�l�Ԁ��!f/�X���"�A������X==[j�`7&�DW�<�4�ֿ�C`ߚ_�錴vi��k��̱��/4Ɨ��^H0 �ҢR8~��Z���"q9gr?4,?>�Z�E��aF.�L� G�ILKo���y3Ju�f9)o�+T�`̊F{�jJ�<|H���C�~jK寂kT�^��<b��}���h�q�^0MrA��<�)����M�@`2����f#�^����¸�$�����$3���:3xZ.}���ͳ�юvM�ƕ.�M-���w+���� d�C��܎�zp�~9Z�e��dR%�E֙5
�D	@9K�eib��｜����'����{e��]-&�R�X�6j8�RƎ��Q����^=M���s��O����"��m�rE���Y�#^pc�h�h��D=Zo���MQ��4��x�A��'o�_>BN�(�:G���0-��߽-�.�뢚_R_�ܝ���z`��9>�Պ����>&U�n�>��(����;�q��-20Pt���x��w9�Z0qN ~��N���u@�7�����Q��<�>��3�f��yHF\w��%Ә(�,o��R,��b�E��)�e �@�5�TB��:ne�B��j`nC��_�q����5�^4��M����GͶ|җ�֧\��'��j�U�2#��%��3�<�;]'O�BL�ڟ�O@+*h�p��II �$�n]9���{�eU.*�O�^9;漬V?K��=�2~��"�����d�RTf1M�����tJ��G�6o����^2D�;��ⷼ���_;u�B�d�s��%D�e� �G�U����t�F����?�˨�'9����΃�S�t���O41���c�<�ڈ�7N
�R����Q�u@S�}��������y���[�:�~�#V
����N�@�lK)f{M�6',p��,_����+�+�ƚ�'G�h���K]�8����(3��j�9�`�_`��ޢ�0�,,�{�<����h2��K�&[}���m����v�s�)���>��?ε,�\Ze�>U{hV.a�B�c~3�� �I����]kXw�Kw4��Z~.�F�t���[���?��ޒ��bC��:_&c1��������M��J�����4&z���^�Geń�x0���\��@0�y�66i�,i��SQ%�r.�子&�p��/o���ר��{G�����s�i���o\�<����\"�˅{Bj,7<�-����h]�B{���C$R�+`>�¶���{ ��8���^��引�K��ׂЭ�ߊ=;"�w��������#���o�d[nu_Qm�Tw����T�*�Z�Y�
F�b��]�l*,�jx����=N<�ѣl��KLQ��SNNR^��<H?}2�UJ�5Y��?�������5��PO<̐}�dS�@g��6��E%���E�q�@��1踠�uFS�	��DϘg����5�r1c|��/;a��1�e�T�x٨�/c[k.��f���U��7b։�3��̏���G�R=���KM�(1�H̺p�b�w͋�����QCn!�d�@O���3h0�x¤�EǠ��&+>�&�Qlr	���Fe���lWa��Lֲ�P��{�>�B\�M��bBrmUD���_����"d�#g�{�q-?Fy���������	�+|D���,�l<�A3q���<���lz����T��X��2~�����f&e��P8Ru8�z7!q+֝M��,�	跼+��gn�^"Ϋ���?�ژm��Z�?��t:,ifp!����`�4�5��A��~�IpRY�߷��j�"��7���������O��;�Ӻ|(L��ė��%���nTS��,CGe'(Pz��)�YK�k���Td媳�ڏ�Y��N������i��wr���~R�ֵ(d0?��_Zs^��9���Y�/uk�q&梁��ż��nv��b�te:�7/�NH��a-l���sssOn��D�`U�8�/M�
1��S���;��#sqE��m��8$���M��G�B_}'���~�a�u�8�iq����I�nG-�{��qttR��7׉6��Z��a�_ �,���+8j��K}�8H���'/��O���}äs��sW/�l�O��5˱�݊�2T3�^U�o��,9bD^�j1W7�������@=H<#X����f����=�"Os*�K�'צ����� �����Oacn<���ṅ��,A�����jq���O�wd_�����7�觿X��"VE/��lufOl`b?D�����酡ܞ˶�����e?�?7 �͒���w}_�E3Mv�Ǹ���i�!��_��/��جt�Wԏ�*y�|OЩ\8�D�[�6o��o��'��B�b�_�:����p��B�nBL��Y�/R`;}W쇹��#1�I���_ѷ�7� _��s5����u��x�CT��B7����#���o��0���2ҽn�t����M+�|.ݽ>LL����h������r�����F��gF2As�-�
��Ʊ%���=�۶����+7+�s� ��M� nЖ���Y 5Yx���7���}�%�y,�b�l?�{����L��d��Gc5����=L�b���h��v3O��L�`��)���;��a/8_�y�\R뼵��_j��tk))LJ��i�{�	�>=*�\���غ[�%������-��(�>���pm�s�0�����%x4�7M����z�����b�2'kĚi�3����7����z"���I��#���d,ҋ'�|��5��D�ZZ�u5�� �{���q܍��Qw=o]�F��^�h����B� �}F�1s�c��ToUlK��^"����^�ǩ�������o���^$2��T�[�#����,nZC`��ѣU���mOE"*�9���wd1&V{����%���Q~T]c��8�Mª�('��=���]A��7��H�.-���������JQ��I���M��QM�"q
�no�X:F?�Q����/��{0��=?��-	\�Ab$YM�V	���^oN�'E��7�g�d��}I��f�������:��I��3Zil���S��\���[ 6�>�]��?���Ay.~�����[�*.i�)����>E�sM=�=�"Ke���gzi����j4�<3����$u��AD|�����j.z3 �#��Kg���8�:��d��{v�C�v�mcF��v2�/�0��˾�1�d~4�2�N;�����el���G�Q��c���r��Ͳ���y�$l��_�)ז=�i�~8�5�
��/�� ���ȦcJ�9�T��w�';����e�ͷ�$!ϵ#צ�9�1��KM"�iN7�YZ�a�V3>���U�mݽ;?C��?�x,,����M����3@�r+=(��;��-LSJ�L���#���7�ۑ6i��I!/��>�Gi/�j*�ҿ����bk�F�n����W������g׫yq��?mrA��T����y��P���rCb0����}Er����5t�9�	�:RD�R�@FL
�W���tA��]j`�sO,���]�F)�A/��]#��bDq�w�>��<B�.�cI���Wu��ݘ��x��ȗ�5��� Ts���%~�p.��eޚ���!��0��]N����^�c����\H�b���p�q�g#넍3���?z5����\�^=� 8D;g}/�x�mf�=zWAy��N��~���3Z%d��Q8ǃ��
�ZV��
t��
�����>������a8mp���]E���_	$��B�AM�^g���E&�10���jW������`~$��<IH�6�l�ٶA��{��_#O��?�#�E�F�8���8'���7f]��A�:'��Q��][�g�ƕ���?��nv&���{�^�x�X*�=� |ʟ�<\K�����_sAH-j�|���N�ֻt�yc�f+�XǸ�CH�]�Xw ��fK�yx]qR��G��φU�Oq��SRGj�>���wV�,g�y,[����w��*���ZI�U�`�K<����K�P�vV�9�TM�U}HY��6���7b%��Fq<��pSͬ��gxw����̞!����w�Z�O[�4��|Ѵ~p�����������}��$��5ȿ������h������Z��C�d�6�\3��z�>�O���٨8A�F��U��&�����ѡ`�J]�&�� 4�$���\�N�zoR�UU�	�Z���I�L*}�5"�x�}�Ӷz��1Li_�ќ����7�HD��P Q$�jv��~��j�pV�L�|{���c ���W�I??��T�ۚ��P-���M�=�O���!\���S��ʛQ���s��0�9� d���ydF1����,&)R�ϻ_\������}���_n4/
>���̖H�t'a����<*O�M,�R��ڲ�Q��8��9���ɐI�"�"���v�¢Oh��8!d��w7��H�0�����.NK�����9*5�0c�rb|�pO�D�AV���6�Wd�LD�Mt�
�ӏ����M}��Jd�P�=i�v�R��<�lu�sﻬ$hdN�K}����:�B0%�<>��/��E�UD-ɥ���������8�5�/�D��Hش������v�e{��{�
'b����j�m�9�~H�8}����*�*-��qR�x�3�.�;[7�<�a�~Y�T'd#�ԑ3m�s߶6'��3U��s?�Ts����e^Q���~w4v1k,�f{ Q�$�����ɏWMG��	���jO�����*���h
Op� f���J*�����r�_�W�(%����q ߪ�7�=|�2�Ӂ{c�rD��t4�YdcF�u�O�0P���(�8w��n^|��3)���Z#2'�5J~
�0<֭t�����V�m���mމGzlI�M3���j�@����`1,b���v���(J6��P/,�댄�a���;L%o9[Ju�d@��%�Ȁo�uI�&s_}y�] ���9d���aTU��9ϥT��>0��Id��j�3��^���&K+>�����"r��J�����l��U�F�7N�֡Z���f��Q �G/�j��c_��N����������s�|ا^��cT����"?�<I�Y�E`��cO��!Ů��2���{�J����E����@w��W�N�1#�:!��
҆'�d���bB�M�f���pY�e6�9��#
i���@^M���-��*�Έ�K!`N�VE���/b�8�B�kj�����֨2��#-�����c��\P��O�h1"�g�~�֤�qөP����NI <3>�p�^@ʹ�3��gt4�=�B9-6���7ٮ�
]��)��j�z8�\�hK-�7�jp[�+��z�����:C�N�fEA�ٴ�q���X�����ܿ]��|�W��wc���T�'{��z[���IG�H���uOU�Cެ^?~�;H�X�X�z�*�e/̌$����Ÿ�E�Qv\�2"���V�F��2e��cK�\D�$�Օ����Mz�Z��l�TdW�B�\ū�e�v��כ��$��yLU����9���(��������5q�̓�+.#PKj8m �I����.v����jЧ� V�@���G$�D�����҄H\��	�Z6��9yN-��l^���]�bG�F�B &��O&b�'����L»�e�kU�L7hhHc����sW�����,��-^���j�����h�uF�'}���f���Q�k��l�wgO��W,����I�a���m�3�&tQ=11ڛ���?@����w���V53o�\� e��5lǥ悏�K��i�tde*�N���T��,~���$nb��;�n#Mw�R}��'D!��7��{V4;�2t�*z:,��@j>�D�a�YI��C��짬�c�;�Q]�Z��%CE��g۩&}��Ǜ&���I��eC�֊��.�N3���h�$C�>F?K�F&�����*�����XY?�>3n|���S�~�s#~�<3��fk���|�m��z�[z�J���b9�a+?���$��V$o|An�y�.��^�ힲ���3��;p1�wp?����G����{�L��X�x4N�u��q4�o�?����Gj�}�t�Np[�<@�[����f�'Y�]AS�C���/c�v�HH�����a"�,�5z$��p�7$��K/����a{����[�V��$iR]X�e���읋P¿��,7�ԕ���ʧm��W&�|.�V������*~!����o̫��o�������ם��S������KW�I}���'�s���JgR�s�f�$�Ӿ�^p9�#?���DR�p���g�g����,�,[��݌�XI���h@�1���o�L�->K�dBkO�c5��^>i���YU^nU��ͪ��s_]�
���I�jh ��S3����mV��k���$:U_\λ�A��m2 9>����h�"_f�Z���H�'�����R{���8��'Pc���W�Yz#8���~��e�����8>�,\����ʒ���c;��J[�K����B��b�cE�|p�X�'k�p,��� �ε�27b2���S��^i�P�m�|�}��� D{����~D����}�f��7h�[2Ǻ����o<V)q9dW:E����,�1��XRi����{�ֈ��%]�?365�$.q��p�ߤ'܁�rd���!�<֛q��>M;��&��?/D_�IJ�"��g���{��\�� ^���U.R�_3|K*t�<"�>Y֕tH.Rs��P��3��[�?�V�1P�b�̚�q�@���OzT	��rH籱�R�0��[���Afoo���(�	*IĤg�놉MS�D�o���ǹ5��[��0[8���J�&�hF�f��Og'��E��I�2Tpio���S��}B�{���|����\/N��Ib����C� �S�0�38::��/:a�k��3kTf�fs*y��Ze
����m�],a�Rr��HV:��_��� ?]ز�����\wI��<y��r������)(<�h�7��lK������'_b~J\�V�y��L�8h;C�Dl�o+Q�'�	��Z{j���¢U��jDm'SN�Э�����K^�:&8�$�\��q�w��+ �k b.06s��|��_�B��_5A
Pi��/�	�ޟ�4�z���sΓ�S\�l|X`�#��ŭ�}RX�_(@um~'�:\_��d'0�+�`a=����� �z\~ٯw�"V_�7����ٞ�JÙ�?(��O���A1�s��e���|߯Ƶ�R�uS���$�r/��@f�Ag'�Ep�ì�A�$��d�|�b�q��|�o��Ywbh>ֲ�[=9e=lh=>�`����z����nD����N��D�
@'6Dձ2���-��?���z��Dv짟�\��G`��b)��wD�>����Z#���Y��$���#'1�VŤ�rɝrb�6�[�ԼnUͦ��a^��z�mg�iȻ`�z�գIMBWq�p�xc�N��5-�j�����7��uj���C9m�Ҿ`�)�~�����T�4t��Ħ������#��V��a��tӍ'����~�+%�mҔ�&���FK4�6O`7���Q��"���J��A-�	p6�ϨaO�R��{�`uK��V�,����t�w^�D�UN�����^tܼ�S�۹G�b9��b��Ղ���|�+�K��?+xs���yr�}va��u�+�([	�k;���l8 ���O�I�+J�j���w|D�{ǪF�:��hU2���*�1�LF1*\�I*��$&��l�m�A��;���j	s��/�o���m��~\�ZmXT;�����-��~4��S�Ac$̗�Ay�>�Yr��ˌ�.K���ջ���\���/�x^3����_���њĝ��7_,�Y������ ֭������)߉��Z����z-v�Z�3.Iq�+j�J@d��nhzl���m�C!sX��`hz⌅/!�̮"7[m�K��Ȯ��Ei!��E߸���B����̀b\v�D"�,�WE�l�D��B?�(���;A�.�%8�`ae1����rc_:hHm��0Fˡ�ݐ��uY��5�f�NͿ2T��5c�M0F�^�~�M3�׆�
�,v��3Z��T��׳���EC���,� ��`z��
�O4�.O������7U�k���6��]��&�n�J����JM_�ϝ�i����6�wm�t}��^�y���>�,n��ɯy�;7���_�9����ɏ�u[��޽o}��)C�	��(p��|�d��`���34�����`���_N����o�������)�	 PK   �|�X��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   �|�Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   �|�X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   �|�X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   �|�X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   �|�XF��-$  ($  /   images/d88a5b0e-66b3-4edb-b452-47f46dd40326.png($�ۉPNG

   IHDR   d   o   %e�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  #�IDATx��}y���/+�ξ�o��[-��I�,�as�k�k{b����Ĭ���X�ځ=�����zc<�'^cds�!�!	��VK�-�}TwuY���<��ZjI�T���̪���z�|��}��p�����>on���,?�aW���Gy瓜{��گg��ש}�w����7@�tvT��2 ]��|j룰dO�f�>�}[)uP)�{���B����ත����0ۂ���G"�[�UEoUѡ
:#N���@l��Ӵ?�(��d6��F"t�"W�� ��b�rR���.(@޼~��`BS��i��b-'N�$�^G���L�&�m#���X�%O;��e��"�>��$<��v']g��/9��ou���	S��;/��!~ d*0I42q�C1q�b)��Jb�:%&�2�J�#=�N )q�Ɖ���]H��U�Oeo}s�����؂�8�ca$2!�>tp� ��.6l�`d��i�,��b��L���dSv%���ޭ�<�[�ʲ��߲JBj
A����c���cy��<����f\C�`MC$&�SI�B�{M�W����}�o*�Q;�й\������u.\�3��f΀V�1?����rȆM>������� �K"��f�⿧8t�R�<[:��ZjtN�H�'�P�N�0�C(�A/��M�6u`�z<'��.jF��R�4R{��8"P���F*�h��R��w�]\G7AO+���rC$�r��;�)��� �q����wl 9���iʠ����0��ފޗ�";���N߃��/C��Q�(�-y/�N=��ڊ��6$��3�f�C_K5�,E��-��Ș�5I���������9C�5���
����)ddK��@(.0����bٗ��Cli=�<�i�������М�pB�B0��;g,��`dd���+uZE��Ɇ���/�=�܃E�!�a6��+���v�F�2�B� #�����l{�3�$�1嘪�H�QT��	WR�@���b��4h�-�|~�, c�0ad0��1Z�@J�Ĥ���0���*!�?���� d�-alղfԮhE�D���C�X\�ٜ0J*���͛��s�!�N��c�Nk�o��F|�K_B�|yfh>��v���}��R�����8Z?N�������]�1����%Ʒ�ёhFk��^W�� �B��r���e�H��5h�$���z�C����L��.�1��O����l`X���9��Ha�PV�ԡ"������J�q�X�|9�|�I������S�r�J|�+_��^t,
A�4y
���0=��a�X��oB*�'a3�t��4P�����XVَ%��D�S#"):�`��I��҇�e� ���J�W��0�8�@�����V"g�W�ƞ�c�=މ��0g���
��3����2X�]�yÕ����y���_��9o�<|�k_�O<����3$�s��8�&����Aqm��݋��QX��.���o܌�<�l���0�e��Oh�ê�K�&�X$��ּ���3�"1�\��LW����A	a�z�P���0�H(���z,�h�����L���Ǯ�Q��aE�*���8�2LDt���>�0�g����P�!444�z���6�7�,,��ߎ_��gȲe����^tQ����_��ub��M�/@�|Ri����`�s-@�D�$���~	��,����#U�0\�pU�H@��[]�� ��baK����*��h�8�f,�h�p�������J��a��}}"�?84g#������O�{<����a�?~����k��/��&&&�Fz�t�k��@����������x�w;j��9�(dl��>�6 �>3����+��v�HG��E_~��H! F�Ĝ�J��n$�¶> aEP�!��v2�`��h�J���wJ�(dD�B����1�t���+�������7����G��v�څC����ڵk=PX}%�I�T���wf�TWW�pVSo�����"��/~��5�nˡm�'ȵ-@0L�=u�`&�^]��hX�d�R~(��,�s���$!�խ�
�3�S���H�-3�� j �WJ@��Q�φ�*�(�l�W%����-�:v@���p
�<��	��_�Ǟ��z6��<ۍ�����7�)��}�Y���<�0����3�<#^ß|�OP���I^��y@��yCGC��5]������dq��h��9�
ny� ���X.(��*O	=�+�5�A0lU�����4r���*ɵ�Ӷ۰���3�o���s�{̠u�i*.{�������-ro�\��c����sp�+=#@�����Ν;1<<�U�yU��8�0����v�G�0�"0\�}y�"|�i�0�??�4��'0E�x�Q��#n�0��3�;��WB�I�FĴ��[1$O[�uqUǥU�yh���%6�>�cAàW��Gn�B�����<����cŊ�<�3d*�7Ŵ���6��a�Z�9W2�@ gmf��WaUr!�I=�D:X%�De�gC�*��|=9�E฀ؒ� ��{�dDD:t�W�ለ-㇤R��+m�`���7���d�\P�.���M0���w�?�B̆f�A_444$�s�Z�䟮��gUe���w����-ע�\���� �f0� J^�q���\Ȏl�-g�*͕���+�tn1+,@��QS}o����VH���/�'Ɵ�.�.����$��,N<�'N�Άf�}2��5���[��E� �i8@����^ppw��� �m�8��D�i�t��������F��)��OM��CgUE@��߆�ߪ�[9�������v���� ��:���C"�\N���Ff0=cw�T� ����~)���<
8�������L��x����'s��dLP�5A�-�XE��.�(�NݿxyF��P�,4�j2\��u܃�s��<9]�iX�������N���K���+�_���Ӌ��-ۀ��z�=�Z�[�RHQ�́���
�D̆l`���U%�����T�׫�*��w�GǞ�Q a���M�����~ؐ��贀�t��u�U��� ��au�6���;Z�̏a���ƀ0X��'q�3���4ޚ�tx�n����I�λOvn�	�
v	GZ�wL�汫uk����销0��k���4J�e�)�Nus
��s���'?}D���p��B#H,%�az�S���T�P��fP�w;���g�!L��`wJ:=�Ćͣh�cA:y��90�+f��k��3�@�QW+�pK�:D԰dL���'Ĉ�b&b5�^�Lh����)��H���[D}��80epD�jߠ��1�p�)�dF@�wmO���Y���p�aUuC�*��jě�S!@X�ݛ�(��խ�S9=KL�p�3��������o@���$}?�OG�5��{gd 1���r����{���K��I:a�����^�ǍX-�������I$;`��Oԯ�k��A��÷'�%>ܘ�Puι��thF@N�PPE���
V[qԺ�~�H����Xe��hy���d����M�s�-7�s�O�@q���5~�B�����`*	H�MKP������n�*k]�R�J�s����V�E93G2ܤ�jؠ4�kpϜk��]/�t��K��J���������= <�u�c���~�?�����X��K4an�A\���<P@�}/��ڙeڎ)i�o=�]�������t,z�l:h6r)V�3� p_B�ĕ߹��]GQ���~�ignY,W&/!�v��k�/&b���?���%CR���Y��tv5_��n��X��n�Q0P�����w]G ��M�������"Z�/Y2���p�y��%��jQ�����XSx���%C2ʦ�Q�TQ{������N�Ԑ��آ��!����}������0^��om@b2'�bZt-��b��C�6N�Z1�c�Q�3>�Ĥk34�����t~�q箆����>v@��cM��n%0���v#��
 �R�Ib��@y�1�:=���(fR"��E���g���n�F�{fM�Z��^��Fv�"E��
���3z�=�u�[yK6K�G�!���n����l�l&7%��b�%6��k��*��"NcЮ�[�w��;���'%��|F	)���S���]˲�.��M��ڽ�q�'P'��K��dGܱer(�0=bp���awK�"%<�rab.���U�SAi�<}|#�V�`�4���>k���=��rs�n�U�t2%ŒG֑[]�wh�îH.�މ�"%��(,WF,|����y/��������@Ϙ�{�"��0��e0J���H_2���&/�l�A�,1�'tM�3q�PH�"��5>@�b�iY�f0g���$t��q
r���w��/[�Շ��(ъm�q�C߸{jk]�M�y*��52u[�t�2�����!�2�̲%$�-6˫:	׽�Y�U��v��r�<��k]C�\pF��1�h�S�H�3����Ɇ���<�I���$�rVY��V$	����<n0�#Gx��L�,�i�`9�@�}�}VcI�!ܑՕ���&��d����I�%D�i��n�9E�R�fG���c; ܑ���T}{���>?��H��w	���"�0P߰��rg��ivda���-�sj�v����r6���i�Aol��Z���*�8�a��r@��G>6E������9R��&@��A�p�?��0E�e<Ό$��p��w�Wk2 �՚�a10�`��,!��l'���g��9sr�(8�܉G,5q5"�VV�;\l�ن4��9,φDH]��P�� �R��?-ϝa̳ȸ�����V��k���~�7�D��}�Ό��?�����߸�IX���VY	ob��gze��Rr`D�NC�����͏4�Z<�> �g�%Xe���`f���#�ʈ�)�c���&��ޔ�}Γ�z�j9�3-��pY4΍�y�E��ס�t��^RgVh�Q/G��F. ţ��Y똚��"����v��t��	.j�,.��%`)���p�p���ʲ�u�dyF�'[Q�}'J�ޥ�5!j\Qrc�K��v�����	�REj���i��H����G�eX΍���݁�3�/�T�:�r~�,�7��R���e��ȭ0��B7W���ኢx.o �n�^V���� ��<��Xٖ��p�p�$��e,�]^#�l�k���P ��UR�I�����(ә�W�v���6�$#���Cp�� QvS3	1A�/�
�rtfs9X?�+��Eq���rE��l���ha5|���6]�Nˎ�,����%C^�M���#;�E_uҫ�ڋ�}���[�~�>$�x�'�dGr���e��®�ŵU҅�r#8J��S;01��ծ��?1��!��PQ':���Dٰ�!KѺ���ftge^M�)�f���ߒ�'�*��{m
��o��Z���a�T5�L�'~��^9(��#Wx8ȳ��!��P[���C~5F1�E�h�6BRR[T팣��Q�
����Rrz�G��%�bi�x���t����i}�`���:5���w����q3�x{h
 r}G2)4U֗��,���I)Zg&5��؝�׮��%t�6����4�;Z��V�g#2u 'R�H�NO�ީ��H��N��WYv@�lH
�������>�p�ŨI�~q$H ;�&IIDbe)9�x�@QMaµ�Lt�e�=�p�@�^�h9sF��^�n��_p`���!Q�rL�|>XA�O*t�����q��R	�D"�T����w��JB�K��PW/����q��W|Ǟ��y���:����p��rQ�1�p�X/:�sexPYJJ�7������T�{o젷�� �����d�a@X�"Z�,��_���5��`N�OG*���;����RR����#'#΅xI��1���C��r8�2�@�� ��+�����<��U=���2���$E�EA	}���	�V7�#�Ĭb0�f�+.�̩�wG�I<�����pq�PH�A׀u��ֈ�*zy?�>����u㪦U�6����waE�b��#�DX��I���g���!��x�����*�����o{���-w���������Mc�
�߆�T`�<Vt��R�ވ�D�<2�!�H��C�V)9+��&	���j*:����ޑ'���Tr���P{C�CRk1Hُ}Gpe�j�{���$.l78���{^���HGXCj_/�~��?>�'w: t
/9�xo�m���(��06����X�Dn�E��g��@$��iU�:�]�~�(��I�izz��>ˊr����[lRާ��D鷺ؖ�ƫ�\U/�.FbV�7�s>�f����,cׅW<��`��ƹc�QpP.0ˊrL8�5���G0n��LYg�.�;(E*"�Ҟp?׹�V���l��m5.�9@H9������kv�W�������*���V�u)6ѳ�qr�h[	�'�_d�0מ���u�*Ĕ^�}GJ��v��Kwb���Zԥ��\r�urn7dcgE7v*��O�/������|��|��o��~��je��<����c�
�R�X�W#|j�������&����G1l�c�r�dO�RإjXټ�c
�6� 6�l3X:~?��&�K��E�ƌbݱᥥ� L<�Ū��7T���<�X��Y(=�'�˚�89��!; �PK`4Fj�-C{�s����;��dQ��s�I�\�]1���-�Z����~� phxpW�,aSB�9!y.���2?F��/ḋ�Ԝh��<��%c���T�Y�ʗ���F������bs
�>1�b��4�]x�C�R�R	���J$	����:V�,�������"��z	7�>�O�ْ��J�!���?oA�Ϸc�ųV��E�[����0�a�����;];��@���H!��*�.,�
���%sۻ�[��]�+��D'���xE�Q������f�^�~�֭�?����f��t.�-];��qړ-�~�T��6���;5��FI #䃡:j�������~~�yw���4s`� g}/��rlܸQL�U�n�m�oh.
ݠa�����\a`8���H������7v%Li3���������U����;gޝ�`A��͙37�|3��y�MN:��> C_t[W�,<r��o�#�,j�@[��p�Զ���x}��F��ؖ�'�llOJ���z`�:
��������/��b�1�k���^:(%�(�wމcǎ�Z�B��?:�Ј����)�l����C�rb��硱�N~��d���Y*x���C�0�O���P����@�v�0lKˑ����E���$�g�%�E�g�9p�@��Č*����C�g?�6o����G��fa�	̸b/�7�i͌a[�.�'j�����I�E6�5�d��uHx=�#c=΍�=ˊ����+q��a�������w��W��_����UW��===3��Lx5�Ç˪�.�|a։_��W�~�zlڴ	������o��1�@��+p<:�ɰ��-����C�aj#Hƫі����zĴ�S�����Z���¸>)����,�7��W��oƉ��,�}�7�ݐ����ר߶m��I���O?��~�e׶�Y��W��������b�вQ�=�W��1I?N�����p��ch��Ese�T%*��.�� r���J�\��A��g�>3��efs��UG�**$�E*�=jq+����3`��I�G^��W���{�`����jۧ�S��,!?��Op���˗���ª�*�	&9F�������W��^�G�i�r
`xe��ѓ�zeKN�05�*�Ǫ#�����a
�(�s�ŒM��Wd�,���[F�᪶j
M5؎�
q�c���yM=�h��g-��F�R��~YY" $}}}��������i������ǽ�ދ�˗#��ʧ^�����F������'7�t:���ڥ)�>��+@������K�;\j0A���iG� �t�	f�((�V�+8�3�lb��Z����.��9��lB@-y��h�0*��$��/��N^b���A�S�b����oK���m��fvww��'��m޼y"-�!^OZ:ɠfm7�EZ�c"=w���ʔg�����fn<����������?�U��^���x��=Ԁ+������.�6� ���=Ś��.E{����Jr�/u2�@ngE/�x���_X���[������d����3p`�l.�ܐ�@_u0�'�E�W'��5M�=��l#x���")��.Y�;{d�=b�b�0^ӂ��s��zժU��v��I�r*L���6���QV�e��Q(��7P��&_��&D9sp<�+S@��P�}E�_WeØ;��5���5X��VX�1��k�=:00�36g��=��r�#S���2z�\�qÆx���H\�zL�
GM\�A_2���8Y�FZɋ�/�2}��ſF������VU	�<$�k����?����9��ʍ���S�ܷ�����{F��݋�I��!gCw�u{�O��L���'�>�@:n�|�ʾ�n���^Gx�1կP�כb�Qϣ
�o�l0��C�dy�	�֦�h�n4�xV�������u�[R�(��y�Gp>�2b�h8]����孧���TkSs|4�ZL��% �Q[APt���=
˗�q f��	��+J'�M�mz[��V�ns���A0CF&�C$H���7� K!�k�b����O�'�qi�%dk�&����S�8 HP;�!���c�" �	�~-��Gҕ�����q��Fs�Y,p�G�&V1R�]�=|��Ge@7�☗l�D>�&�H�`�sK��� /v�W�^�0�� �}��*�q���$H/�������G� ��[w�������B����l �(�G�������&��@�b�    IEND�B`�PK   �|�X��6�B  �  /   images/ea05fd3c-afe5-4b36-b101-0986c4cae35e.png��s���b``���p	�) ��$MR,鎾����$�����L�K@�Q]�S:PP��5�$%�$�*�(H1Z�X���X�[���[�ʞ͊�!7?%3����f�;X�<]C*漝�!�*q�����x~μ��}Ukk�Ƭ��W6���z��ɸtU|] �2U���"��y,�N�K�,��\2)��掛o��w[o~�y�M�L͊�����hom�y�̟o���3'VOן{��7�S�S&O�Y���I�i��N�~����
}��'+�?I�>���q�f��l3��4o��W,?*-o-�p���!�2Dh�S�3���O���sO���gΡ���G P�o����%�2_Ż��9�=��tiȱ?A����j{<��Y�����������g�ZT����}��ձ·�+�l��?-a�1��u}���ˮ�2a���K[��n�5[�w�3ެ��������!��4��˷L���LN���7G�=n�+��L!=�~����J�R�3m��/�r�E�5�SVs��KGj�����ҷ�O��_���8�7���@��G
E̒;���g�+�(z�{z��ݒ!^�w]�p�z��[���;W��;�c���)B��.��V����X�ua��̕72���j�?��U��U\u6Wms��Ό�:�͜皻x]꒢��+�:�v;kѦ]<WVE�k��k�.g�6a���,��ཻZ��Y�ND{���-��L�&-7�U��}���V{���[]��X�wئ�C����i�Vw����?u�=fs���I��ji뱴���9.;�u���Dq�
ߕ���:^����Ֆ%��ڋ�D{��=�r睯�褷��{��d�sL����<|�����^1��`��G�)��f���^"z���m�Ov)�]��x5�1*xꭐ.��/gO>�DGƲ�C��G锧�dL��������jx�Kc��r
m��`~�W59鉿'\V��^���yw�Xu-\t{Ҫy;�d�K%����]qv��̲u����¬�ݽI[�K�?Xx�[�4����s��]�ݹa�������ST��&�Iը���n��ޛ;�ٿ��]�m�@��@,�*m�����t���5���*���h��F�M����V��w��X<*�b��Z��5�c�~�}W��L��|�bV^5ܿ����[������,���~����X��&����|��u��+��e];������i}�1+3��,�ҥ%?Z6=��Y�J��e{<wfH���Y�@���hJS�����_���+N?{��������Y�����u=sG��W���{��6}r�.�jΏ���,w�[x�"��e�t�sY�� PK   �|�X�T�|  �  /   images/f1ab8fe3-f826-4bea-bba4-7763291602bf.png�YyPSY����m@��\XTFа	0:bЀ
e5��	�@�D�a\�d0C"F� aT`�.a�$*;�D� YH�e���x��^��W5��ֹ��>}������.:;~�}�v��ܙ� І��{����O�h6�;�@��������s�Q ���3$��N�@�'@��� �9�7�EͥS�����π����Y�@�-����ƣ/���{��N0��	<�u�nK0Q{�8��y��-zh���g�A0/�&��{�%�V�;:�
M�/?���n�ߥ��h�4f�ݙB��N�,�B�g�}��|�}�u`Ka1:�N����7Q�g����{�-��&�}�^>(�X5ݾ9��O�1'E*��ź��i�1�2�B���ԒK��!C��>��߹K��G����>F?���شAN���B���6��K��q������_L�4��2ǲR�R�A����ii�A�m�^D����<�.�.>���Xz�$v�xZ�d�
�"l9f�ŔTڀ�$�4�⦾T:�v�,5�#��I::�� Y�GuaA��-����c�}�1��Ū��E4E��B������KR�c}�g�yzm����Ly*H�5��4��4vH}�����Χ�g���m�ߤ7�
&+ΐڒ+����H�ZwIc���T�G��L�*�P,F.��#0`���I��J%O1��&׏��٧-�΅H>�N֙lp�T="w4���s\��V,����5\z����O?�Mv���� �_^؄˂Hl��2M�T�CfG}��rN`(������uc�����f�\���.�8-�ᵒ�(p���h^���	�x4��i�5/!12^���y�n��b�\�;� Ev/��E�̹����P�~��+բH��8z�
_�ʞXD֯|�+�{��3��O�)�G1\��sԵB�X#�/��/4����<x;<�v��b���n��J���9�H���M��j����8���:<��e�*��s�K6V7'k�Ԇ�,w�;�V���N��C�Qg��h���s�_�%�Iڝ��V=�N�b#�1,��X@�Het��������]haK���S.��.�uCu:�>Z�ʳkwq=WXs� gū�hY�"�&�[�$(Қu�;Ӝf��Ē��� Fy���>��-�;���r�x�P��#��.��%qqrU��|4���N)�s-��s~����ȡ��SUvP��P�w��C�J���w/��u���wDM��`¡:}����ǀ���(ٷ%�CC��{,JL��Uʘ�<�Kl��R6�m�x�Shl����5V��.�m�O:��f��i���gPU��U����˩�匝r5��%�'=/	9R�4��:{S��]pV? �񕤃��>���,PQ����#o@����~ ��yT�Z3Ev������=3s���	�-�[�0O�7E�������~�Pƻ��7T#����o��jd���}��W�d�\^`>/ī����3}���:1�Օ�`�sQdhN�0����l�u� z�Ý��z���b'�)K�lcș{�ͻ�#ws��7l�m?0�r �ݸ�ξkC.��d���/K��M��D�ґk���ԯ��o@���Z3���:�k^��J�_TZ�D�@��C��jiE��6Qf��,�`�b�Hw��O 9LB�ă␨�y���S_XF�l�Km\�tԌE����:�r9���һzyM�N՝Pu~��<t�<=�1x:����e.V�X_�6�̖`e�g�-��do�e���J�B������<#�Id��U��ٛ�d#&Z9:��Ӭ𥧧��"!S����P�E�k�~=Gtɵ�\R��5.9F�h�˛���JGK�o�Ɣ�1?�,Qe���g����o>���ޮ�h��s��`��6d�j�d�L��=�Swt)�R%Gx1�k_S��?:#b�j��#�J/H��ٞ$�/��xtqKKc��1�s|}	���)���ɾ���*�S��[���|�.�<R��y��N_�9?�(g/J�E�
�����5��,'"f�Ci�rJ��v9N�D���b�rd���ʶ��G�twJo�$n�2�eᝧH�7�1��]�Hz��whʋ���#�ָؚ!�CQ��_�'J��.i�U���#/�b[h���c �����#KQ\����|'�6�Iy{Z�~Ь���ݝ���=�AM:dX���?�Y�����m05�����,�������M��+rI8�:���;��V��0Jxj~�i#�z0�/B��o�����#�� ﺛ �y��k�Tr8;%�����\9�;ZJ��>�P2��ޥӻ���2C�ya���rϓ�l#t�.�����I~��yt�e��E�C�ݼ+.����Ւcf��03@���NT)����R	�^��Q�в��O��)2}2_Sʊ��cb7��Oޫ
J��+�M3�}{�v^�����]9y��mK#ca�Z���]�.�W���՝��q����6?b��KgA`���&��Y�Վ
��#���>뽿X�JFey�c��!��Ex��/^��j����.���K#����E��Z:�B�������IV1�ΐ���˹���Y�3���΁c���E) `�МO[�ʿ�˺y�c�Bb���=�9H8���u*�����?�yG��Đ��O����f>�J������N�u�rGmtȧ�CE�X�:U�F��%�Z-�[O_���Io{��47 �U�Ћ�ƣ�G���m���gj.W߹r�* ��$gƃ]��k���w�^Rqvng&��4���ͩnW�C��}=1�݉�х��|������z�;n��+Y/W�^G~�˝�vu��Q#2�Aز0d�	w1ֵ\�h�h(4�V�7�k����/e�տy����G��h"j%5|�TP`���$�vg�p�3��|�~�`�!�Ym!*n����]�	����g�%�@�EV2��S��?uUc[w���@�Nf��!�n���r�ӱF�N��N�y�w֟�Sޤc��!?�0���Ȓ,P�sQ*W9:��@���&��[��U&�!��msSx�z|q�A@��yW�ٸ3�o���cБR�UtіU?/zfZ�[k��Ý�V��ci{�����ۊ�}W�~܍7\=�7k�P����C��Ĕ�;��t�%XX$�8���:T�dj=|�T��?�Q�cp���6{e�k�w9 �U��ftQI_w.Bf<`1���LU��d�r:V?ܪ*W����Q�,�42��\�������Ks���������>э �
 ��L��k���zVì��x��<�h"
�˛�	�|]\�1�&�&l������o�З[P>�:��Ѥ�_@m����߳|4�޽�����!�����p��o���Ft}��bi<@�p}�� �p�j�b��<�5�U@��kp�����k��;Ԃ�ʋu�F/6y�{����|�����V�����L�Kf=�����6*O`��w�(.6$�/�j���z5�.��ĭH2--��g�L��e���TY��T��!���ٜ�j0����ǚ�ҙ.%�s���p���c��A8�~���=��-݃���^�7��?�T�-��^��hmt5����ۉ"_S��"�ђ�v[z;�����ƗW�/2���&�pj6�'�o��7eo~++ʼp��/(P��뎦���G�diJq�	��J���Iۯ�3@�
CQ��T��SyH�&[5R��E1��'�[y���Go�q�e�Pa﫞����e�a�!L0w�~w�%����}��	֎U^�R�O����-M����u4L�'����p�ل��M4���>r�E� j�/�5|��6ދkQ--=\=�Rѹ����u�M}�G7���a� ���8�,eAll?�[���Q��͗��᝚�]QN4�n�Z���j��zտs�L/@4-�5x4/�-l�sm㾬����]��S~�Ŷ�C�`�}(�����W�M6�M^f�x����J�ie�P���8A���[oW6�E�cKg����13�tIkŅ�+��X�_q=�� �c�u�S̳W�'y�vU&��_2׷��L��8��]A��"�S8S�z�{wa�t�2��g���<F:Ȝ�" fQ�/	pM����Tb��~lK���eb����˺D���/�q"W�����=<�ԍP�Q ���3ן6�f�dR7��*��0xAQ�c��q�8�+$n�3��!T��m�{��I9�����?���t$��M ��8��:�&��n|T_���/�5G�#��#�_��������,\V��Q��ȳ�W��d,Gù�����Y���G�'4f�b_����K�uܚ?�-�3��8���0kj��{d,Ȋv\�f=��ar�ǻs�,��E�^��9h�^[���J��,��8a�򇍒1u�'��-&�RK�8m��u�U�f� !��-�eY�Q�<Kܛ�����
{�i�{��53�zܖuG�ߟ3E�P�0�[_h�W�6�LZ�l f���(�����H�!����IJh�QJ���K����
�]���+ksfR�6�ג��F4)��r��z����z���<�^6�Я���k����C��!��4Ź2˙��֯d�Z:��{�x��%̷5V3w�vb"��D�����]G��o����s��$�H�q�$�����?$J�7���µ����רy<�;O̪7T���A�w�O�'�O�z���#�{$�9�LY5!�o����g��B8�(�T[����q�bz��;}�F�!���Ĕ�C�K�7ܽtWn�)�2�n�p~�=���t�`[c6�]d�Qi�)�Gu<���v�+ec���1(��2+���yܬ6�
��{	\j���
�/�3�gV�XM}��WJ����V7Cv�o�����H����<:�������qŗ�=��i�P����ı��X��D)�����FW�ھ,z�s����_�x`�gE^�;i"��r��n�k�&>����]�Ƚ���h����@���/�7�u�v�g�R3[>D{w�k�(i��(}5>+�q��'�R���~�7���̊��[�B�PZ98.,���ɢ��/����`��qY$�/� jPT��,�͛��FJ�ࠂҬ��\䂋>"�K��5������hi��4�Į.�("�aM��^^*���ϱ��ʂ ݉�m���n��Kl�e����uHzHTx������]|`��uR�Ĝ֥y醤Tu�X%@9.F�:�+��Xs�KȜ���{��	���92!��a_��35g;Z0b�ܬ/��i���*C�6V�+<I���e�����ߜ�����1AwLfF1�?��´�$��Ձ�9��Mk�"��C oXK|>�n@��l�I5`S�����Ic���T��hꩨ��`Q��I�4)u��_�I
o��j�L�,�x��[�$c���i>���Km��\~L� :��QS�f����i��X q��'��k���	��o��n��NR��5��f���_�e��Z��n^U����ҋ$}��Z�Y�2�'�]X`�(٪튖�n�{	�c��>�"ŝ��f���(���K?*M�	���=��G6�=\�t�٘4B5����M7�{�~�F���ա�{��VG�z�n�&[���Qcl}���'�/�I�4��'���$g3QĴ��B-�u�!�i���G�~�q^�&�%��S�Su���K$Ɯj�54.��������߂a�or�����OX��8�4���?��8A�em�o�C�~1��������ȟ�ϔ�x��PK   �|�X
���J  
     jsons/user_defined.json�X�n�F�A@���/~K�5��HܼF0kLT&U.5#ԟ�7����I��Th^����9�sϽgt3m�,��h�ֱ�bʋ���_���8��;u�W���Ǜ��{Ս�x���e�O��&'��.f�<�K�/��HELב G�FJE�=1֋��S^-�"͇5:�ɭ�;j�6��9����E��zG�,�f�G@��'�c�Ȅ���
sTb�e��3��}Y,G	�#�E����QI�b�8��zЕ�_���K�9��?y�/�OY��i����ʹh�N�z1�_��y�1#P�^�{�����LR��r�.����r���
��nU�"VMޯ�����eyE;y�4��Wp#L��ʷy�-Ѓ�&;��j�(�NE��"�WBN���M�(��%v��b$b�N����D�E���@2j��ԥU\�Fn� d�p��f�n�w3m���h��}S�yݽP�y��u>�;H@�w�L�Ϻ5�����`�:����n��ºy���v�߆BFP��j�0�Ţm&d��`�1޶�8�;����dp~>2?;��bd~�_��W[����V{C���n������ӧu�	0�If`?I�a�m��~�&FP6�M*
�)mzPU�MY�o�F�7�F]��l*��+�UAg3X���fm��%$��e��Z�c���~��ͪ^��o�c06��]����9��ޫ�m߸�.�}��-�d}�V�����u�2Σo���}} ���"��Ȧ(��3	���Bd"�:���#�vi�}yyr49�.'�R�����#N�w+��A#� �DB�08�:��p��%���}?���!���n����h��"ۙ�`V>������[5g�V�L�.m�6a��8ɴyҬ�W_�!�:�-\ ������<��-z2��\F�Tx�5��#����N��xG�����bJ���Uih��J��0lSBDF�ڒ*d�6H�pBK��Գ��tmӔ�#u�_����{m\t�;�HY.P`ʡȈ���D�u��S��'�V���O�'��P�N�#��c{�U�S����0���w����af�d�^���Ͼ�n~�`�;�}v�3��Pd/�Ꮍ�=��\��m�}yj�c58{w�H��t�N.��š�A��
�#��1PEp�qAW��8fT��O^�MY��i�J�38ŀ��i`���y�IL!y�ݮ� ��1F�D�q�(yk���R�ӭ��z��$fFmk����3E#��_�js�W�2a��z�����4�X�m���Lj���j�´9h�V������`S����m7&�YŵI��Bx
����(�X0:N8�B��:�7���@f�{��ࢅ �o-Cz)����Չs�;��g%���$w`G�f�I&�7�"��t-�m��?
�e����vqC�{Kt7*{o\�ʀD�j���P���[�,��>ީ�ٵ&����*�q{(�~d���3��g�n_ܓg 2��.���y��N�3�(���HCy��-�����?�ݟ�%~�%���M6o�+���4ya�P�q�	�ɝ�Tͼ�&D����Ѝ��!˘ XQn��Q~T��GE8@E���/PK
   �|�X�IyQ#  %^                  cirkitFile.jsonPK
   �|�XWC��)�  � /             ~#  images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK
   5^�X�ZD) �, /             ��  images/1b210ea0-4cba-494f-997a-67bd7381b5cc.pngPK
   5^�X:u�� �� /             �! images/3d480ee1-e9cf-4ef6-9de8-5a7043d7f31b.pngPK
   �|�X'(�5W �@ /             Y� images/4737cce6-ef6b-4e79-82eb-dab57378d86e.pngPK
   �|�X��_8
  3
  /             �� images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK
   �|�Xd��  �   /             �� images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   �|�X?S��� 2� /             �� images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   �|�X	��#u } /             |� images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   �|�X$�8�l  �  /             �K images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   �|�XF��-$  ($  /             �i images/d88a5b0e-66b3-4edb-b452-47f46dd40326.pngPK
   �|�X��6�B  �  /             � images/ea05fd3c-afe5-4b36-b101-0986c4cae35e.pngPK
   �|�X�T�|  �  /             �� images/f1ab8fe3-f826-4bea-bba4-7763291602bf.pngPK
   �|�X
���J  
               � jsons/user_defined.jsonPK      �  ��   